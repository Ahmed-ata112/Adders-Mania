/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Nov  4 15:00:36 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3015833075 */

module CLA_4bit__0_47(a, b, cin, sum, cout);
   input [3:0]a;
   input [3:0]b;
   input cin;
   output [3:0]sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;

   AOI21_X1 i_0_0 (.A(n_0_11), .B1(n_0_10), .B2(n_0_2), .ZN(cout));
   XOR2_X1 i_0_1 (.A(b[0]), .B(a[0]), .Z(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_6), .B(n_0_0), .ZN(sum[1]));
   XOR2_X1 i_0_3 (.A(b[1]), .B(a[1]), .Z(n_0_0));
   XNOR2_X1 i_0_4 (.A(n_0_5), .B(n_0_1), .ZN(sum[2]));
   XNOR2_X1 i_0_5 (.A(b[2]), .B(a[2]), .ZN(n_0_1));
   XNOR2_X1 i_0_6 (.A(n_0_9), .B(n_0_2), .ZN(sum[3]));
   OAI21_X1 i_0_7 (.A(n_0_3), .B1(a[2]), .B2(b[2]), .ZN(n_0_2));
   INV_X1 i_0_8 (.A(n_0_4), .ZN(n_0_3));
   AOI21_X1 i_0_9 (.A(n_0_5), .B1(a[2]), .B2(b[2]), .ZN(n_0_4));
   OAI21_X1 i_0_10 (.A(n_0_7), .B1(n_0_8), .B2(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_11 (.A1(b[0]), .A2(a[0]), .ZN(n_0_6));
   NAND2_X1 i_0_12 (.A1(b[1]), .A2(a[1]), .ZN(n_0_7));
   NOR2_X1 i_0_13 (.A1(b[1]), .A2(a[1]), .ZN(n_0_8));
   XOR2_X1 i_0_14 (.A(b[3]), .B(a[3]), .Z(n_0_9));
   NAND2_X1 i_0_15 (.A1(b[3]), .A2(a[3]), .ZN(n_0_10));
   NOR2_X1 i_0_16 (.A1(b[3]), .A2(a[3]), .ZN(n_0_11));
endmodule

module CLA_4bit__0_63(a, b, cin, sum, cout);
   input [3:0]a;
   input [3:0]b;
   input cin;
   output [3:0]sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   OAI21_X1 i_0_0 (.A(n_0_1), .B1(n_0_2), .B2(n_0_0), .ZN(cout));
   XOR2_X1 i_0_1 (.A(cin), .B(n_0_9), .Z(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_8), .B(n_0_6), .ZN(sum[1]));
   XNOR2_X1 i_0_3 (.A(n_0_5), .B(n_0_3), .ZN(sum[2]));
   XOR2_X1 i_0_4 (.A(n_0_2), .B(n_0_0), .Z(sum[3]));
   OAI21_X1 i_0_5 (.A(n_0_1), .B1(b[3]), .B2(a[3]), .ZN(n_0_0));
   NAND2_X1 i_0_6 (.A1(b[3]), .A2(a[3]), .ZN(n_0_1));
   AOI22_X1 i_0_7 (.A1(b[2]), .A2(a[2]), .B1(n_0_4), .B2(n_0_3), .ZN(n_0_2));
   XOR2_X1 i_0_8 (.A(b[2]), .B(a[2]), .Z(n_0_3));
   INV_X1 i_0_9 (.A(n_0_5), .ZN(n_0_4));
   AOI22_X1 i_0_10 (.A1(b[1]), .A2(a[1]), .B1(n_0_7), .B2(n_0_6), .ZN(n_0_5));
   XOR2_X1 i_0_11 (.A(b[1]), .B(a[1]), .Z(n_0_6));
   INV_X1 i_0_12 (.A(n_0_8), .ZN(n_0_7));
   AOI22_X1 i_0_13 (.A1(b[0]), .A2(a[0]), .B1(cin), .B2(n_0_9), .ZN(n_0_8));
   XOR2_X1 i_0_14 (.A(b[0]), .B(a[0]), .Z(n_0_9));
endmodule

module CLA_4bit__0_71(a, b, cin, sum, cout);
   input [3:0]a;
   input [3:0]b;
   input cin;
   output [3:0]sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   OAI21_X1 i_0_0 (.A(n_0_1), .B1(n_0_2), .B2(n_0_0), .ZN(cout));
   XOR2_X1 i_0_1 (.A(cin), .B(n_0_9), .Z(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_8), .B(n_0_6), .ZN(sum[1]));
   XNOR2_X1 i_0_3 (.A(n_0_5), .B(n_0_3), .ZN(sum[2]));
   XOR2_X1 i_0_4 (.A(n_0_2), .B(n_0_0), .Z(sum[3]));
   OAI21_X1 i_0_5 (.A(n_0_1), .B1(b[3]), .B2(a[3]), .ZN(n_0_0));
   NAND2_X1 i_0_6 (.A1(b[3]), .A2(a[3]), .ZN(n_0_1));
   AOI22_X1 i_0_7 (.A1(b[2]), .A2(a[2]), .B1(n_0_4), .B2(n_0_3), .ZN(n_0_2));
   XOR2_X1 i_0_8 (.A(b[2]), .B(a[2]), .Z(n_0_3));
   INV_X1 i_0_9 (.A(n_0_5), .ZN(n_0_4));
   AOI22_X1 i_0_10 (.A1(b[1]), .A2(a[1]), .B1(n_0_7), .B2(n_0_6), .ZN(n_0_5));
   XOR2_X1 i_0_11 (.A(b[1]), .B(a[1]), .Z(n_0_6));
   INV_X1 i_0_12 (.A(n_0_8), .ZN(n_0_7));
   AOI22_X1 i_0_13 (.A1(b[0]), .A2(a[0]), .B1(cin), .B2(n_0_9), .ZN(n_0_8));
   XOR2_X1 i_0_14 (.A(b[0]), .B(a[0]), .Z(n_0_9));
endmodule

module CLA_4bit__0_79(a, b, cin, sum, cout);
   input [3:0]a;
   input [3:0]b;
   input cin;
   output [3:0]sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   OAI21_X1 i_0_0 (.A(n_0_1), .B1(n_0_2), .B2(n_0_0), .ZN(cout));
   XOR2_X1 i_0_1 (.A(cin), .B(n_0_9), .Z(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_8), .B(n_0_6), .ZN(sum[1]));
   XNOR2_X1 i_0_3 (.A(n_0_5), .B(n_0_3), .ZN(sum[2]));
   XOR2_X1 i_0_4 (.A(n_0_2), .B(n_0_0), .Z(sum[3]));
   OAI21_X1 i_0_5 (.A(n_0_1), .B1(b[3]), .B2(a[3]), .ZN(n_0_0));
   NAND2_X1 i_0_6 (.A1(b[3]), .A2(a[3]), .ZN(n_0_1));
   AOI22_X1 i_0_7 (.A1(b[2]), .A2(a[2]), .B1(n_0_4), .B2(n_0_3), .ZN(n_0_2));
   XOR2_X1 i_0_8 (.A(b[2]), .B(a[2]), .Z(n_0_3));
   INV_X1 i_0_9 (.A(n_0_5), .ZN(n_0_4));
   AOI22_X1 i_0_10 (.A1(b[1]), .A2(a[1]), .B1(n_0_7), .B2(n_0_6), .ZN(n_0_5));
   XOR2_X1 i_0_11 (.A(b[1]), .B(a[1]), .Z(n_0_6));
   INV_X1 i_0_12 (.A(n_0_8), .ZN(n_0_7));
   AOI22_X1 i_0_13 (.A1(b[0]), .A2(a[0]), .B1(cin), .B2(n_0_9), .ZN(n_0_8));
   XOR2_X1 i_0_14 (.A(b[0]), .B(a[0]), .Z(n_0_9));
endmodule

module CLA_4bit__0_87(a, b, cin, sum, cout);
   input [3:0]a;
   input [3:0]b;
   input cin;
   output [3:0]sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   OAI21_X1 i_0_0 (.A(n_0_1), .B1(n_0_2), .B2(n_0_0), .ZN(cout));
   XOR2_X1 i_0_1 (.A(cin), .B(n_0_9), .Z(sum[0]));
   XNOR2_X1 i_0_2 (.A(n_0_8), .B(n_0_6), .ZN(sum[1]));
   XNOR2_X1 i_0_3 (.A(n_0_5), .B(n_0_3), .ZN(sum[2]));
   XOR2_X1 i_0_4 (.A(n_0_2), .B(n_0_0), .Z(sum[3]));
   OAI21_X1 i_0_5 (.A(n_0_1), .B1(b[3]), .B2(a[3]), .ZN(n_0_0));
   NAND2_X1 i_0_6 (.A1(b[3]), .A2(a[3]), .ZN(n_0_1));
   AOI22_X1 i_0_7 (.A1(b[2]), .A2(a[2]), .B1(n_0_4), .B2(n_0_3), .ZN(n_0_2));
   XOR2_X1 i_0_8 (.A(b[2]), .B(a[2]), .Z(n_0_3));
   INV_X1 i_0_9 (.A(n_0_5), .ZN(n_0_4));
   AOI22_X1 i_0_10 (.A1(b[1]), .A2(a[1]), .B1(n_0_7), .B2(n_0_6), .ZN(n_0_5));
   XOR2_X1 i_0_11 (.A(b[1]), .B(a[1]), .Z(n_0_6));
   INV_X1 i_0_12 (.A(n_0_8), .ZN(n_0_7));
   AOI22_X1 i_0_13 (.A1(b[0]), .A2(a[0]), .B1(cin), .B2(n_0_9), .ZN(n_0_8));
   XOR2_X1 i_0_14 (.A(b[0]), .B(a[0]), .Z(n_0_9));
endmodule

module CLA_4bit__0_95(a, b, cin, sum, cout);
   input [3:0]a;
   input [3:0]b;
   input cin;
   output [3:0]sum;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;

   XNOR2_X1 i_0_0 (.A(b[0]), .B(n_0_0), .ZN(sum[0]));
   XNOR2_X1 i_0_1 (.A(a[0]), .B(cin), .ZN(n_0_0));
   XNOR2_X1 i_0_2 (.A(n_0_9), .B(n_0_1), .ZN(sum[1]));
   XOR2_X1 i_0_3 (.A(b[1]), .B(a[1]), .Z(n_0_1));
   XNOR2_X1 i_0_4 (.A(n_0_7), .B(n_0_2), .ZN(sum[2]));
   XOR2_X1 i_0_5 (.A(b[2]), .B(a[2]), .Z(n_0_2));
   NOR2_X1 i_0_6 (.A1(cout), .A2(n_0_3), .ZN(sum[3]));
   NOR2_X1 i_0_7 (.A1(a[3]), .A2(n_0_4), .ZN(n_0_3));
   AND2_X1 i_0_8 (.A1(a[3]), .A2(n_0_4), .ZN(cout));
   OAI21_X1 i_0_9 (.A(n_0_5), .B1(n_0_7), .B2(n_0_6), .ZN(n_0_4));
   NAND2_X1 i_0_10 (.A1(b[2]), .A2(a[2]), .ZN(n_0_5));
   NOR2_X1 i_0_11 (.A1(b[2]), .A2(a[2]), .ZN(n_0_6));
   OAI21_X1 i_0_12 (.A(n_0_8), .B1(a[1]), .B2(b[1]), .ZN(n_0_7));
   NAND2_X1 i_0_13 (.A1(n_0_12), .A2(n_0_9), .ZN(n_0_8));
   OAI21_X1 i_0_14 (.A(n_0_10), .B1(cin), .B2(a[0]), .ZN(n_0_9));
   INV_X1 i_0_15 (.A(n_0_11), .ZN(n_0_10));
   AOI21_X1 i_0_16 (.A(b[0]), .B1(a[0]), .B2(cin), .ZN(n_0_11));
   NAND2_X1 i_0_17 (.A1(b[1]), .A2(a[1]), .ZN(n_0_12));
endmodule

module CLA_4bit(a, b, cin, sum, cout);
   input [3:0]a;
   input [3:0]b;
   input cin;
   output [3:0]sum;
   output cout;

   XOR2_X1 i_0_0 (.A(a[3]), .B(cin), .Z(sum[0]));
endmodule

module CLA(in1, in2, cin, sum, cout, of);
   input [31:0]in1;
   input [31:0]in2;
   input cin;
   output [31:0]sum;
   output cout;
   output of;

   wire c;

   CLA_4bit__0_47 cla1 (.a({in1[3], in1[2], in1[1], in1[0]}), .b({in2[3], in2[2], 
      in2[1], in2[0]}), .cin(), .sum({sum[3], sum[2], sum[1], sum[0]}), .cout(c));
   CLA_4bit__0_63 genblk1_4_cla (.a({in1[7], in1[6], in1[5], in1[4]}), .b({
      in2[7], in2[6], in2[5], in2[4]}), .cin(c), .sum({sum[7], sum[6], sum[5], 
      sum[4]}), .cout(n_0));
   CLA_4bit__0_71 genblk1_8_cla (.a({in1[11], in1[10], in1[9], in1[8]}), 
      .b({in2[11], in2[10], in2[9], in2[8]}), .cin(n_0), .sum({sum[11], sum[10], 
      sum[9], sum[8]}), .cout(n_1));
   CLA_4bit__0_79 genblk1_12_cla (.a({in1[15], in1[14], in1[13], in1[12]}), 
      .b({in2[15], in2[14], in2[13], in2[12]}), .cin(n_1), .sum({sum[15], 
      sum[14], sum[13], sum[12]}), .cout(n_2));
   CLA_4bit__0_87 genblk1_16_cla (.a({in1[19], in1[18], in1[17], in1[16]}), 
      .b({in2[19], in2[18], in2[17], in2[16]}), .cin(n_2), .sum({sum[19], 
      sum[18], sum[17], sum[16]}), .cout(n_3));
   CLA_4bit__0_95 genblk1_20_cla (.a({in1[23], in1[22], in1[21], in1[20]}), 
      .b({uc_0, in2[22], in2[21], in2[20]}), .cin(n_3), .sum({sum[23], sum[22], 
      sum[21], sum[20]}), .cout(n_4));
   CLA_4bit genblk1_24_cla (.a({in1[31], uc_1, uc_2, uc_3}), .b(), .cin(n_4), 
      .sum({uc_4, uc_5, uc_6, sum[24]}), .cout());
endmodule

module count_leading_zeros(valueIn, result);
   input [22:0]valueIn;
   output [4:0]result;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;

   AOI21_X1 i_0_0 (.A(valueIn[22]), .B1(n_0_40), .B2(n_0_0), .ZN(result[0]));
   OAI21_X1 i_0_1 (.A(n_0_39), .B1(valueIn[19]), .B2(n_0_1), .ZN(n_0_0));
   AOI21_X1 i_0_2 (.A(valueIn[18]), .B1(n_0_38), .B2(n_0_2), .ZN(n_0_1));
   OAI21_X1 i_0_3 (.A(n_0_37), .B1(valueIn[15]), .B2(n_0_3), .ZN(n_0_2));
   AOI21_X1 i_0_4 (.A(valueIn[14]), .B1(n_0_36), .B2(n_0_4), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(n_0_35), .B1(valueIn[11]), .B2(n_0_5), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(valueIn[10]), .B1(n_0_34), .B2(n_0_6), .ZN(n_0_5));
   OAI21_X1 i_0_7 (.A(n_0_33), .B1(valueIn[7]), .B2(n_0_7), .ZN(n_0_6));
   AOI21_X1 i_0_8 (.A(valueIn[6]), .B1(n_0_32), .B2(n_0_8), .ZN(n_0_7));
   OAI21_X1 i_0_9 (.A(n_0_31), .B1(valueIn[3]), .B2(n_0_9), .ZN(n_0_8));
   AOI21_X1 i_0_10 (.A(valueIn[2]), .B1(n_0_30), .B2(valueIn[0]), .ZN(n_0_9));
   NOR3_X1 i_0_11 (.A1(valueIn[22]), .A2(valueIn[21]), .A3(n_0_10), .ZN(
      result[1]));
   NOR3_X1 i_0_12 (.A1(valueIn[20]), .A2(valueIn[19]), .A3(n_0_11), .ZN(n_0_10));
   NOR3_X1 i_0_13 (.A1(valueIn[18]), .A2(valueIn[17]), .A3(n_0_12), .ZN(n_0_11));
   NOR3_X1 i_0_14 (.A1(valueIn[16]), .A2(valueIn[15]), .A3(n_0_13), .ZN(n_0_12));
   NOR3_X1 i_0_15 (.A1(valueIn[14]), .A2(valueIn[13]), .A3(n_0_14), .ZN(n_0_13));
   AOI211_X1 i_0_16 (.A(valueIn[12]), .B(valueIn[11]), .C1(n_0_15), .C2(n_0_25), 
      .ZN(n_0_14));
   OAI21_X1 i_0_17 (.A(n_0_24), .B1(n_0_16), .B2(n_0_21), .ZN(n_0_15));
   NOR3_X1 i_0_18 (.A1(valueIn[4]), .A2(valueIn[3]), .A3(n_0_17), .ZN(n_0_16));
   NOR2_X1 i_0_19 (.A1(valueIn[2]), .A2(valueIn[1]), .ZN(n_0_17));
   AND2_X1 i_0_20 (.A1(n_0_18), .A2(n_0_29), .ZN(result[2]));
   NAND2_X1 i_0_21 (.A1(n_0_19), .A2(n_0_28), .ZN(n_0_18));
   OAI21_X1 i_0_22 (.A(n_0_26), .B1(n_0_20), .B2(n_0_23), .ZN(n_0_19));
   NOR3_X1 i_0_23 (.A1(n_0_21), .A2(valueIn[3]), .A3(valueIn[4]), .ZN(n_0_20));
   OR2_X1 i_0_24 (.A1(valueIn[6]), .A2(valueIn[5]), .ZN(n_0_21));
   AND3_X1 i_0_25 (.A1(n_0_22), .A2(n_0_28), .A3(n_0_29), .ZN(result[3]));
   NOR2_X1 i_0_26 (.A1(n_0_27), .A2(n_0_22), .ZN(result[4]));
   NAND3_X1 i_0_27 (.A1(n_0_26), .A2(n_0_25), .A3(n_0_24), .ZN(n_0_22));
   NAND2_X1 i_0_28 (.A1(n_0_25), .A2(n_0_24), .ZN(n_0_23));
   NOR2_X1 i_0_29 (.A1(valueIn[8]), .A2(valueIn[7]), .ZN(n_0_24));
   NOR2_X1 i_0_30 (.A1(valueIn[10]), .A2(valueIn[9]), .ZN(n_0_25));
   NOR4_X1 i_0_31 (.A1(valueIn[14]), .A2(valueIn[13]), .A3(valueIn[12]), 
      .A4(valueIn[11]), .ZN(n_0_26));
   NAND2_X1 i_0_32 (.A1(n_0_29), .A2(n_0_28), .ZN(n_0_27));
   NOR4_X1 i_0_33 (.A1(valueIn[18]), .A2(valueIn[17]), .A3(valueIn[16]), 
      .A4(valueIn[15]), .ZN(n_0_28));
   NOR4_X1 i_0_34 (.A1(valueIn[22]), .A2(valueIn[21]), .A3(valueIn[20]), 
      .A4(valueIn[19]), .ZN(n_0_29));
   INV_X1 i_0_35 (.A(valueIn[1]), .ZN(n_0_30));
   INV_X1 i_0_36 (.A(valueIn[4]), .ZN(n_0_31));
   INV_X1 i_0_37 (.A(valueIn[5]), .ZN(n_0_32));
   INV_X1 i_0_38 (.A(valueIn[8]), .ZN(n_0_33));
   INV_X1 i_0_39 (.A(valueIn[9]), .ZN(n_0_34));
   INV_X1 i_0_40 (.A(valueIn[12]), .ZN(n_0_35));
   INV_X1 i_0_41 (.A(valueIn[13]), .ZN(n_0_36));
   INV_X1 i_0_42 (.A(valueIn[16]), .ZN(n_0_37));
   INV_X1 i_0_43 (.A(valueIn[17]), .ZN(n_0_38));
   INV_X1 i_0_44 (.A(valueIn[20]), .ZN(n_0_39));
   INV_X1 i_0_45 (.A(valueIn[21]), .ZN(n_0_40));
endmodule

module datapath__0_28(p_0, p_1);
   input [4:0]p_0;
   output [15:0]p_1;

   INV_X1 i_0 (.A(p_0[1]), .ZN(p_1[1]));
   INV_X1 i_1 (.A(p_0[2]), .ZN(p_1[2]));
   INV_X1 i_2 (.A(p_0[3]), .ZN(p_1[3]));
   INV_X1 i_3 (.A(p_0[4]), .ZN(p_1[4]));
   INV_X1 i_4 (.A(p_0[0]), .ZN(p_1[8]));
endmodule

module datapath__0_30(p_0, exp_Sum, exp_Sum1);
   input [15:0]p_0;
   input [7:0]exp_Sum;
   output [7:0]exp_Sum1;

   FA_X1 i_0 (.A(p_0[0]), .B(exp_Sum[0]), .CI(p_0[8]), .CO(n_0), .S(exp_Sum1[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(exp_Sum[1]), .CI(n_0), .CO(n_1), .S(exp_Sum1[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(exp_Sum[2]), .CI(n_1), .CO(n_2), .S(exp_Sum1[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(exp_Sum[3]), .CI(n_2), .CO(n_3), .S(exp_Sum1[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(exp_Sum[4]), .CI(n_3), .CO(n_4), .S(exp_Sum1[4]));
   FA_X1 i_5 (.A(p_0[7]), .B(exp_Sum[5]), .CI(n_4), .CO(n_5), .S(exp_Sum1[5]));
   FA_X1 i_6 (.A(p_0[7]), .B(exp_Sum[6]), .CI(n_5), .CO(n_6), .S(exp_Sum1[6]));
   XNOR2_X1 i_7 (.A(p_0[7]), .B(exp_Sum[7]), .ZN(n_7));
   XNOR2_X1 i_8 (.A(n_7), .B(n_6), .ZN(exp_Sum1[7]));
endmodule

module datapath__0_37(p_0, p_1);
   input [23:0]p_0;
   output [31:0]p_1;

   XOR2_X1 i_0 (.A(p_0[1]), .B(p_0[0]), .Z(p_1[1]));
   AND2_X1 i_1 (.A1(n_21), .A2(n_0), .ZN(p_1[2]));
   OAI21_X1 i_2 (.A(p_0[2]), .B1(p_0[1]), .B2(p_0[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(p_0[3]), .B(n_21), .Z(p_1[3]));
   XOR2_X1 i_4 (.A(p_0[4]), .B(n_20), .Z(p_1[4]));
   XOR2_X1 i_5 (.A(p_0[5]), .B(n_19), .Z(p_1[5]));
   AND2_X1 i_6 (.A1(n_18), .A2(n_1), .ZN(p_1[6]));
   OAI21_X1 i_7 (.A(p_0[6]), .B1(n_19), .B2(p_0[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(p_0[7]), .B(n_18), .Z(p_1[7]));
   XOR2_X1 i_9 (.A(p_0[8]), .B(n_17), .Z(p_1[8]));
   AND2_X1 i_10 (.A1(n_16), .A2(n_2), .ZN(p_1[9]));
   OAI21_X1 i_11 (.A(p_0[9]), .B1(n_17), .B2(p_0[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(p_0[10]), .B(n_16), .Z(p_1[10]));
   XNOR2_X1 i_13 (.A(p_0[11]), .B(n_15), .ZN(p_1[11]));
   XOR2_X1 i_14 (.A(p_0[12]), .B(n_14), .Z(p_1[12]));
   XOR2_X1 i_15 (.A(p_0[13]), .B(n_13), .Z(p_1[13]));
   XNOR2_X1 i_16 (.A(p_0[14]), .B(n_12), .ZN(p_1[14]));
   XNOR2_X1 i_17 (.A(p_0[15]), .B(n_11), .ZN(p_1[15]));
   XOR2_X1 i_18 (.A(p_0[16]), .B(n_10), .Z(p_1[16]));
   XOR2_X1 i_19 (.A(p_0[17]), .B(n_9), .Z(p_1[17]));
   XOR2_X1 i_20 (.A(p_0[18]), .B(n_8), .Z(p_1[18]));
   AND2_X1 i_21 (.A1(n_7), .A2(n_3), .ZN(p_1[19]));
   OAI21_X1 i_22 (.A(p_0[19]), .B1(n_8), .B2(p_0[18]), .ZN(n_3));
   XOR2_X1 i_23 (.A(p_0[20]), .B(n_7), .Z(p_1[20]));
   AND2_X1 i_24 (.A1(n_6), .A2(n_4), .ZN(p_1[21]));
   OAI21_X1 i_25 (.A(p_0[21]), .B1(n_7), .B2(p_0[20]), .ZN(n_4));
   XOR2_X1 i_26 (.A(p_0[22]), .B(n_6), .Z(p_1[22]));
   AND2_X1 i_27 (.A1(p_1[31]), .A2(n_5), .ZN(p_1[23]));
   OAI21_X1 i_28 (.A(p_0[23]), .B1(n_6), .B2(p_0[22]), .ZN(n_5));
   OR3_X1 i_29 (.A1(n_6), .A2(p_0[22]), .A3(p_0[23]), .ZN(p_1[31]));
   OR3_X1 i_30 (.A1(n_7), .A2(p_0[20]), .A3(p_0[21]), .ZN(n_6));
   OR3_X1 i_31 (.A1(n_8), .A2(p_0[18]), .A3(p_0[19]), .ZN(n_7));
   OR2_X1 i_32 (.A1(n_9), .A2(p_0[17]), .ZN(n_8));
   OR2_X1 i_33 (.A1(n_10), .A2(p_0[16]), .ZN(n_9));
   NAND2_X1 i_34 (.A1(n_11), .A2(n_23), .ZN(n_10));
   NOR3_X1 i_35 (.A1(n_13), .A2(p_0[13]), .A3(p_0[14]), .ZN(n_11));
   NOR2_X1 i_36 (.A1(n_13), .A2(p_0[13]), .ZN(n_12));
   OR2_X1 i_37 (.A1(n_14), .A2(p_0[12]), .ZN(n_13));
   NAND2_X1 i_38 (.A1(n_15), .A2(n_22), .ZN(n_14));
   NOR2_X1 i_39 (.A1(n_16), .A2(p_0[10]), .ZN(n_15));
   OR3_X1 i_40 (.A1(n_17), .A2(p_0[8]), .A3(p_0[9]), .ZN(n_16));
   OR2_X1 i_41 (.A1(n_18), .A2(p_0[7]), .ZN(n_17));
   OR3_X1 i_42 (.A1(n_19), .A2(p_0[5]), .A3(p_0[6]), .ZN(n_18));
   OR2_X1 i_43 (.A1(n_20), .A2(p_0[4]), .ZN(n_19));
   OR2_X1 i_44 (.A1(n_21), .A2(p_0[3]), .ZN(n_20));
   OR3_X1 i_45 (.A1(p_0[2]), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_21));
   INV_X1 i_46 (.A(p_0[11]), .ZN(n_22));
   INV_X1 i_47 (.A(p_0[15]), .ZN(n_23));
endmodule

module fp_adder(A, B, Sum, overflow, underflow);
   input [31:0]A;
   input [31:0]B;
   output [31:0]Sum;
   output overflow;
   output underflow;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire [4:0]num_leading_zeros;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_58;
   wire n_0_0_0;
   wire n_0_59;
   wire n_0_0_1;
   wire n_0_60;
   wire n_0_0_2;
   wire [31:0]mant_A_reg;
   wire n_0_54;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_55;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_56;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_62;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_63;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_64;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_65;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_66;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_67;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_68;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_69;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_70;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_71;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_72;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_74;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_75;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_76;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_77;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_78;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_79;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_80;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_81;
   wire n_0_0_117;
   wire n_0_82;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_83;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_84;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_85;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_86;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_87;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_88;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_89;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_90;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_91;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_92;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_93;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_94;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_95;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_96;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_97;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_98;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_99;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_100;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_101;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_102;
   wire n_0_0_230;
   wire n_0_0_231;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_103;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_104;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_0_246;
   wire n_0_105;
   wire n_0_0_247;
   wire n_0_0_248;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_0_253;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_112;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_113;
   wire n_0_0_282;
   wire n_0_114;
   wire n_0_0_283;
   wire n_0_115;
   wire n_0_0_284;
   wire n_0_116;
   wire n_0_0_285;
   wire n_0_117;
   wire n_0_0_286;
   wire n_0_118;
   wire n_0_0_287;
   wire n_0_119;
   wire n_0_0_288;
   wire n_0_120;
   wire n_0_0_289;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_0_304;
   wire n_0_0_305;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_0_311;
   wire n_0_0_312;
   wire n_0_0_313;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_0_321;
   wire n_0_0_322;
   wire n_0_0_323;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_328;
   wire n_0_0_329;
   wire n_0_0_330;
   wire n_0_0_331;
   wire n_0_0_332;
   wire n_0_0_333;
   wire n_0_0_334;
   wire n_0_0_335;
   wire n_0_0_336;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_341;
   wire n_0_0_342;
   wire n_0_0_343;
   wire n_0_0_344;
   wire n_0_0_345;
   wire n_0_0_346;
   wire n_0_0_347;
   wire n_0_0_348;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_351;
   wire n_0_0_352;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_0_355;
   wire n_0_0_356;
   wire n_0_0_357;
   wire n_0_0_358;
   wire n_0_0_359;
   wire n_0_0_360;
   wire n_0_0_361;
   wire n_0_0_362;
   wire n_0_0_363;
   wire n_0_0_364;
   wire n_0_0_365;
   wire n_0_0_366;
   wire n_0_0_367;
   wire n_0_0_368;
   wire n_0_0_369;
   wire n_0_0_370;
   wire n_0_0_371;
   wire n_0_0_372;
   wire n_0_0_373;
   wire n_0_0_374;
   wire n_0_0_375;
   wire n_0_0_376;
   wire n_0_0_377;
   wire n_0_0_378;
   wire n_0_0_379;
   wire n_0_0_380;
   wire n_0_0_381;
   wire n_0_0_382;
   wire n_0_0_383;
   wire n_0_0_384;
   wire n_0_0_385;
   wire n_0_0_386;
   wire n_0_0_387;
   wire n_0_0_388;
   wire n_0_0_389;
   wire n_0_0_390;
   wire n_0_0_391;
   wire n_0_0_392;
   wire n_0_0_393;
   wire n_0_0_394;
   wire n_0_0_395;
   wire n_0_0_396;
   wire n_0_0_397;
   wire n_0_0_398;
   wire n_0_0_399;
   wire n_0_0_400;
   wire n_0_0_401;
   wire n_0_0_402;
   wire n_0_106;
   wire n_0_0_403;
   wire n_0_111;
   wire n_0_0_404;
   wire n_0_0_405;
   wire n_0_0_406;
   wire n_0_0_407;
   wire n_0_0_408;
   wire n_0_0_409;
   wire n_0_0_410;
   wire n_0_0_411;
   wire n_0_0_412;
   wire n_0_0_413;
   wire n_0_0_414;
   wire n_0_0_415;
   wire n_0_0_416;
   wire n_0_0_417;
   wire n_0_0_418;
   wire n_0_0_419;
   wire n_0_0_420;
   wire n_0_0_421;
   wire n_0_0_422;
   wire n_0_0_423;
   wire n_0_0_424;
   wire n_0_0_425;
   wire n_0_0_426;
   wire n_0_0_427;
   wire n_0_0_428;
   wire n_0_0_429;
   wire n_0_0_430;
   wire n_0_0_431;
   wire n_0_0_432;
   wire n_0_0_433;
   wire n_0_0_434;
   wire n_0_0_435;
   wire n_0_0_436;
   wire n_0_61;
   wire n_0_0_437;
   wire n_0_0_438;
   wire n_0_57;
   wire n_0_0_439;
   wire n_0_0_440;
   wire n_0_0_441;
   wire n_0_0_442;
   wire n_0_0_443;
   wire n_0_0_444;
   wire n_0_0_445;
   wire n_0_0_446;
   wire n_0_0_447;
   wire n_0_0_448;
   wire n_0_0_449;
   wire n_0_0_450;
   wire n_0_0_451;
   wire n_0_0_452;
   wire n_0_0_453;
   wire n_0_0_454;
   wire n_0_0_455;
   wire n_0_0_456;
   wire n_0_0_457;
   wire n_0_0_458;
   wire n_0_0_459;
   wire n_0_0_460;
   wire n_0_0_461;
   wire n_0_0_462;

   CLA CLA_dut (.in1({mant_A_reg[31], uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, 
      mant_A_reg[23], mant_A_reg[22], mant_A_reg[21], mant_A_reg[20], 
      mant_A_reg[19], mant_A_reg[18], mant_A_reg[17], mant_A_reg[16], 
      mant_A_reg[15], mant_A_reg[14], mant_A_reg[13], mant_A_reg[12], 
      mant_A_reg[11], mant_A_reg[10], mant_A_reg[9], mant_A_reg[8], 
      mant_A_reg[7], mant_A_reg[6], mant_A_reg[5], mant_A_reg[4], mant_A_reg[3], 
      mant_A_reg[2], mant_A_reg[1], n_0_54}), .in2({uc_7, uc_8, uc_9, uc_10, 
      uc_11, uc_12, uc_13, uc_14, uc_15, n_0_105, n_0_104, n_0_103, n_0_102, 
      n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, n_0_93, 
      n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, 
      n_0_83}), .cin(), .sum({uc_16, uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0}), .cout(), .of());
   count_leading_zeros count_leading_zeros_instance (.valueIn({n_0_22, n_0_21, 
      n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, 
      n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, 
      n_0_1, n_0_0}), .result(num_leading_zeros));
   datapath__0_28 i_0_11 (.p_0({n_0_61, n_0_60, n_0_59, n_0_58, n_0_57}), 
      .p_1({uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29, n_0_29, uc_30, 
      uc_31, uc_32, n_0_28, n_0_27, n_0_26, n_0_25, uc_33}));
   datapath__0_30 i_0_13 (.p_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      n_0_112, n_0_111, uc_34, uc_35, n_0_110, n_0_109, n_0_108, n_0_107, 
      n_0_106}), .exp_Sum({n_0_120, n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, 
      n_0_114, n_0_113}), .exp_Sum1({Sum[30], Sum[29], Sum[28], Sum[27], Sum[26], 
      Sum[25], Sum[24], Sum[23]}));
   datapath__0_37 i_0_20 (.p_0({n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, 
      n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, 
      n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, n_0_56, n_0_55, n_0_54}), 
      .p_1({n_0_53, uc_36, uc_37, uc_38, uc_39, uc_40, uc_41, uc_42, n_0_52, 
      n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, 
      n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, 
      n_0_33, n_0_32, n_0_31, n_0_30, uc_43}));
   HA_X1 i_0_0_0 (.A(num_leading_zeros[1]), .B(num_leading_zeros[0]), .CO(
      n_0_0_0), .S(n_0_58));
   HA_X1 i_0_0_1 (.A(num_leading_zeros[2]), .B(n_0_0_0), .CO(n_0_0_1), .S(n_0_59));
   HA_X1 i_0_0_2 (.A(num_leading_zeros[3]), .B(n_0_0_1), .CO(n_0_0_2), .S(n_0_60));
   MUX2_X1 i_0_0_3 (.A(n_0_30), .B(n_0_55), .S(n_0_0_408), .Z(mant_A_reg[1]));
   MUX2_X1 i_0_0_4 (.A(n_0_31), .B(n_0_56), .S(n_0_0_408), .Z(mant_A_reg[2]));
   MUX2_X1 i_0_0_5 (.A(n_0_32), .B(n_0_62), .S(n_0_0_408), .Z(mant_A_reg[3]));
   MUX2_X1 i_0_0_6 (.A(n_0_33), .B(n_0_63), .S(n_0_0_408), .Z(mant_A_reg[4]));
   MUX2_X1 i_0_0_7 (.A(n_0_34), .B(n_0_64), .S(n_0_0_408), .Z(mant_A_reg[5]));
   MUX2_X1 i_0_0_8 (.A(n_0_35), .B(n_0_65), .S(n_0_0_408), .Z(mant_A_reg[6]));
   MUX2_X1 i_0_0_9 (.A(n_0_36), .B(n_0_66), .S(n_0_0_408), .Z(mant_A_reg[7]));
   MUX2_X1 i_0_0_10 (.A(n_0_37), .B(n_0_67), .S(n_0_0_408), .Z(mant_A_reg[8]));
   MUX2_X1 i_0_0_11 (.A(n_0_38), .B(n_0_68), .S(n_0_0_408), .Z(mant_A_reg[9]));
   MUX2_X1 i_0_0_12 (.A(n_0_39), .B(n_0_69), .S(n_0_0_408), .Z(mant_A_reg[10]));
   MUX2_X1 i_0_0_13 (.A(n_0_40), .B(n_0_70), .S(n_0_0_408), .Z(mant_A_reg[11]));
   MUX2_X1 i_0_0_14 (.A(n_0_41), .B(n_0_71), .S(n_0_0_408), .Z(mant_A_reg[12]));
   MUX2_X1 i_0_0_15 (.A(n_0_42), .B(n_0_72), .S(n_0_0_408), .Z(mant_A_reg[13]));
   MUX2_X1 i_0_0_16 (.A(n_0_43), .B(n_0_73), .S(n_0_0_408), .Z(mant_A_reg[14]));
   MUX2_X1 i_0_0_17 (.A(n_0_44), .B(n_0_74), .S(n_0_0_408), .Z(mant_A_reg[15]));
   MUX2_X1 i_0_0_18 (.A(n_0_45), .B(n_0_75), .S(n_0_0_408), .Z(mant_A_reg[16]));
   MUX2_X1 i_0_0_19 (.A(n_0_46), .B(n_0_76), .S(n_0_0_408), .Z(mant_A_reg[17]));
   MUX2_X1 i_0_0_20 (.A(n_0_47), .B(n_0_77), .S(n_0_0_408), .Z(mant_A_reg[18]));
   MUX2_X1 i_0_0_21 (.A(n_0_48), .B(n_0_78), .S(n_0_0_408), .Z(mant_A_reg[19]));
   MUX2_X1 i_0_0_22 (.A(n_0_49), .B(n_0_79), .S(n_0_0_408), .Z(mant_A_reg[20]));
   MUX2_X1 i_0_0_23 (.A(n_0_50), .B(n_0_80), .S(n_0_0_408), .Z(mant_A_reg[21]));
   MUX2_X1 i_0_0_24 (.A(n_0_51), .B(n_0_81), .S(n_0_0_408), .Z(mant_A_reg[22]));
   MUX2_X1 i_0_0_25 (.A(n_0_52), .B(n_0_82), .S(n_0_0_408), .Z(mant_A_reg[23]));
   AND2_X1 i_0_0_26 (.A1(n_0_0_407), .A2(n_0_53), .ZN(mant_A_reg[31]));
   OAI221_X1 i_0_0_27 (.A(n_0_0_3), .B1(n_0_0_4), .B2(n_0_0_100), .C1(n_0_0_101), 
      .C2(n_0_0_7), .ZN(n_0_54));
   NAND2_X1 i_0_0_28 (.A1(A[0]), .A2(n_0_0_458), .ZN(n_0_0_3));
   OAI21_X1 i_0_0_29 (.A(n_0_0_5), .B1(n_0_0_15), .B2(n_0_0_125), .ZN(n_0_0_4));
   OAI211_X1 i_0_0_30 (.A(n_0_0_6), .B(n_0_0_125), .C1(n_0_0_462), .C2(n_0_0_28), 
      .ZN(n_0_0_5));
   AOI222_X1 i_0_0_31 (.A1(A[0]), .A2(n_0_0_119), .B1(n_0_0_73), .B2(A[8]), 
      .C1(A[16]), .C2(n_0_0_22), .ZN(n_0_0_6));
   OAI221_X1 i_0_0_32 (.A(n_0_0_11), .B1(n_0_0_7), .B2(n_0_0_100), .C1(n_0_0_12), 
      .C2(n_0_0_101), .ZN(n_0_55));
   OAI21_X1 i_0_0_33 (.A(n_0_0_10), .B1(n_0_0_8), .B2(n_0_0_126), .ZN(n_0_0_7));
   OAI21_X1 i_0_0_34 (.A(n_0_0_9), .B1(n_0_0_33), .B2(n_0_0_462), .ZN(n_0_0_8));
   AOI222_X1 i_0_0_35 (.A1(A[1]), .A2(n_0_0_119), .B1(n_0_0_73), .B2(A[9]), 
      .C1(A[17]), .C2(n_0_0_22), .ZN(n_0_0_9));
   NAND2_X1 i_0_0_36 (.A1(n_0_0_19), .A2(n_0_0_126), .ZN(n_0_0_10));
   NAND2_X1 i_0_0_37 (.A1(A[1]), .A2(n_0_0_458), .ZN(n_0_0_11));
   OAI221_X1 i_0_0_38 (.A(n_0_0_17), .B1(n_0_0_12), .B2(n_0_0_100), .C1(n_0_0_18), 
      .C2(n_0_0_101), .ZN(n_0_56));
   INV_X1 i_0_0_39 (.A(n_0_0_13), .ZN(n_0_0_12));
   AOI21_X1 i_0_0_40 (.A(n_0_0_14), .B1(n_0_0_26), .B2(n_0_0_126), .ZN(n_0_0_13));
   NOR2_X1 i_0_0_41 (.A1(n_0_0_126), .A2(n_0_0_15), .ZN(n_0_0_14));
   OAI21_X1 i_0_0_42 (.A(n_0_0_16), .B1(n_0_0_41), .B2(n_0_0_462), .ZN(n_0_0_15));
   AOI222_X1 i_0_0_43 (.A1(A[2]), .A2(n_0_0_119), .B1(n_0_0_73), .B2(A[10]), 
      .C1(A[18]), .C2(n_0_0_22), .ZN(n_0_0_16));
   NAND2_X1 i_0_0_44 (.A1(A[2]), .A2(n_0_0_458), .ZN(n_0_0_17));
   OAI221_X1 i_0_0_45 (.A(n_0_0_23), .B1(n_0_0_24), .B2(n_0_0_101), .C1(n_0_0_18), 
      .C2(n_0_0_100), .ZN(n_0_62));
   MUX2_X1 i_0_0_46 (.A(n_0_0_19), .B(n_0_0_31), .S(n_0_0_126), .Z(n_0_0_18));
   AOI221_X1 i_0_0_47 (.A(n_0_0_20), .B1(n_0_0_47), .B2(n_0_0_124), .C1(A[11]), 
      .C2(n_0_0_73), .ZN(n_0_0_19));
   INV_X1 i_0_0_48 (.A(n_0_0_21), .ZN(n_0_0_20));
   AOI22_X1 i_0_0_49 (.A1(A[3]), .A2(n_0_0_119), .B1(n_0_0_22), .B2(A[19]), 
      .ZN(n_0_0_21));
   NOR3_X1 i_0_0_50 (.A1(n_0_0_123), .A2(n_0_0_121), .A3(n_0_0_124), .ZN(
      n_0_0_22));
   NAND2_X1 i_0_0_51 (.A1(A[3]), .A2(n_0_0_458), .ZN(n_0_0_23));
   OAI221_X1 i_0_0_52 (.A(n_0_0_29), .B1(n_0_0_24), .B2(n_0_0_100), .C1(n_0_0_30), 
      .C2(n_0_0_101), .ZN(n_0_63));
   OAI21_X1 i_0_0_53 (.A(n_0_0_25), .B1(n_0_0_38), .B2(n_0_0_125), .ZN(n_0_0_24));
   NAND2_X1 i_0_0_54 (.A1(n_0_0_125), .A2(n_0_0_26), .ZN(n_0_0_25));
   AOI221_X1 i_0_0_55 (.A(n_0_0_27), .B1(n_0_0_96), .B2(A[8]), .C1(A[16]), 
      .C2(n_0_0_51), .ZN(n_0_0_26));
   NOR2_X1 i_0_0_56 (.A1(n_0_0_124), .A2(n_0_0_28), .ZN(n_0_0_27));
   AOI222_X1 i_0_0_57 (.A1(A[4]), .A2(n_0_0_120), .B1(n_0_0_84), .B2(A[12]), 
      .C1(A[20]), .C2(n_0_0_42), .ZN(n_0_0_28));
   NAND2_X1 i_0_0_58 (.A1(A[4]), .A2(n_0_0_458), .ZN(n_0_0_29));
   OAI221_X1 i_0_0_59 (.A(n_0_0_34), .B1(n_0_0_35), .B2(n_0_0_101), .C1(
      n_0_0_100), .C2(n_0_0_30), .ZN(n_0_64));
   MUX2_X1 i_0_0_60 (.A(n_0_0_45), .B(n_0_0_31), .S(n_0_0_125), .Z(n_0_0_30));
   AOI221_X1 i_0_0_61 (.A(n_0_0_32), .B1(n_0_0_96), .B2(A[9]), .C1(A[17]), 
      .C2(n_0_0_51), .ZN(n_0_0_31));
   NOR2_X1 i_0_0_62 (.A1(n_0_0_124), .A2(n_0_0_33), .ZN(n_0_0_32));
   AOI222_X1 i_0_0_63 (.A1(A[5]), .A2(n_0_0_120), .B1(n_0_0_84), .B2(A[13]), 
      .C1(A[21]), .C2(n_0_0_42), .ZN(n_0_0_33));
   NAND2_X1 i_0_0_64 (.A1(A[5]), .A2(n_0_0_458), .ZN(n_0_0_34));
   OAI221_X1 i_0_0_65 (.A(n_0_0_43), .B1(n_0_0_101), .B2(n_0_0_44), .C1(n_0_0_35), 
      .C2(n_0_0_100), .ZN(n_0_65));
   INV_X1 i_0_0_66 (.A(n_0_0_36), .ZN(n_0_0_35));
   OAI21_X1 i_0_0_67 (.A(n_0_0_37), .B1(n_0_0_50), .B2(n_0_0_125), .ZN(n_0_0_36));
   NAND2_X1 i_0_0_68 (.A1(n_0_0_38), .A2(n_0_0_125), .ZN(n_0_0_37));
   INV_X1 i_0_0_69 (.A(n_0_0_39), .ZN(n_0_0_38));
   AOI221_X1 i_0_0_70 (.A(n_0_0_40), .B1(n_0_0_96), .B2(A[10]), .C1(A[18]), 
      .C2(n_0_0_51), .ZN(n_0_0_39));
   NOR2_X1 i_0_0_71 (.A1(n_0_0_124), .A2(n_0_0_41), .ZN(n_0_0_40));
   AOI222_X1 i_0_0_72 (.A1(A[6]), .A2(n_0_0_120), .B1(n_0_0_84), .B2(A[14]), 
      .C1(A[22]), .C2(n_0_0_42), .ZN(n_0_0_41));
   NOR2_X1 i_0_0_73 (.A1(n_0_0_123), .A2(n_0_0_121), .ZN(n_0_0_42));
   NAND2_X1 i_0_0_74 (.A1(A[6]), .A2(n_0_0_458), .ZN(n_0_0_43));
   OAI221_X1 i_0_0_75 (.A(n_0_0_48), .B1(n_0_0_44), .B2(n_0_0_100), .C1(n_0_0_49), 
      .C2(n_0_0_101), .ZN(n_0_66));
   MUX2_X1 i_0_0_76 (.A(n_0_0_45), .B(n_0_0_56), .S(n_0_0_126), .Z(n_0_0_44));
   OAI21_X1 i_0_0_77 (.A(n_0_0_46), .B1(n_0_0_47), .B2(n_0_0_124), .ZN(n_0_0_45));
   NAND2_X1 i_0_0_78 (.A1(n_0_0_124), .A2(n_0_0_64), .ZN(n_0_0_46));
   AOI22_X1 i_0_0_79 (.A1(n_0_0_439), .A2(n_0_0_120), .B1(n_0_0_83), .B2(
      n_0_0_121), .ZN(n_0_0_47));
   NAND2_X1 i_0_0_80 (.A1(A[7]), .A2(n_0_0_458), .ZN(n_0_0_48));
   OAI221_X1 i_0_0_81 (.A(n_0_0_54), .B1(n_0_0_101), .B2(n_0_0_55), .C1(n_0_0_49), 
      .C2(n_0_0_100), .ZN(n_0_67));
   MUX2_X1 i_0_0_82 (.A(n_0_0_50), .B(n_0_0_59), .S(n_0_0_126), .Z(n_0_0_49));
   AOI221_X1 i_0_0_83 (.A(n_0_0_52), .B1(n_0_0_51), .B2(A[20]), .C1(A[16]), 
      .C2(n_0_0_73), .ZN(n_0_0_50));
   AND2_X1 i_0_0_84 (.A1(n_0_0_124), .A2(n_0_0_84), .ZN(n_0_0_51));
   INV_X1 i_0_0_85 (.A(n_0_0_53), .ZN(n_0_0_52));
   AOI22_X1 i_0_0_86 (.A1(A[8]), .A2(n_0_0_119), .B1(n_0_0_96), .B2(A[12]), 
      .ZN(n_0_0_53));
   NAND2_X1 i_0_0_87 (.A1(A[8]), .A2(n_0_0_458), .ZN(n_0_0_54));
   OAI221_X1 i_0_0_88 (.A(n_0_0_57), .B1(n_0_0_55), .B2(n_0_0_100), .C1(n_0_0_58), 
      .C2(n_0_0_101), .ZN(n_0_68));
   MUX2_X1 i_0_0_89 (.A(n_0_0_56), .B(n_0_0_63), .S(n_0_0_126), .Z(n_0_0_55));
   AOI222_X1 i_0_0_90 (.A1(A[9]), .A2(n_0_0_119), .B1(n_0_0_96), .B2(A[13]), 
      .C1(n_0_0_84), .C2(n_0_0_92), .ZN(n_0_0_56));
   NAND2_X1 i_0_0_91 (.A1(A[9]), .A2(n_0_0_458), .ZN(n_0_0_57));
   OAI221_X1 i_0_0_92 (.A(n_0_0_61), .B1(n_0_0_101), .B2(n_0_0_62), .C1(n_0_0_58), 
      .C2(n_0_0_100), .ZN(n_0_69));
   MUX2_X1 i_0_0_93 (.A(n_0_0_69), .B(n_0_0_59), .S(n_0_0_125), .Z(n_0_0_58));
   AOI221_X1 i_0_0_94 (.A(n_0_0_60), .B1(n_0_0_119), .B2(A[10]), .C1(A[18]), 
      .C2(n_0_0_73), .ZN(n_0_0_59));
   NOR2_X1 i_0_0_95 (.A1(n_0_0_462), .A2(n_0_0_77), .ZN(n_0_0_60));
   NAND2_X1 i_0_0_96 (.A1(A[10]), .A2(n_0_0_458), .ZN(n_0_0_61));
   OAI221_X1 i_0_0_97 (.A(n_0_0_65), .B1(n_0_0_62), .B2(n_0_0_100), .C1(n_0_0_67), 
      .C2(n_0_0_101), .ZN(n_0_70));
   MUX2_X1 i_0_0_98 (.A(n_0_0_63), .B(n_0_0_72), .S(n_0_0_126), .Z(n_0_0_62));
   MUX2_X1 i_0_0_99 (.A(n_0_0_82), .B(n_0_0_64), .S(n_0_0_462), .Z(n_0_0_63));
   AOI22_X1 i_0_0_100 (.A1(A[11]), .A2(n_0_0_120), .B1(n_0_0_84), .B2(A[19]), 
      .ZN(n_0_0_64));
   NAND2_X1 i_0_0_101 (.A1(A[11]), .A2(n_0_0_458), .ZN(n_0_0_65));
   OAI221_X1 i_0_0_102 (.A(n_0_0_66), .B1(n_0_0_67), .B2(n_0_0_100), .C1(
      n_0_0_101), .C2(n_0_0_71), .ZN(n_0_71));
   NAND2_X1 i_0_0_103 (.A1(A[12]), .A2(n_0_0_458), .ZN(n_0_0_66));
   MUX2_X1 i_0_0_104 (.A(n_0_0_68), .B(n_0_0_69), .S(n_0_0_125), .Z(n_0_0_67));
   AOI21_X1 i_0_0_105 (.A(n_0_0_76), .B1(n_0_0_96), .B2(A[18]), .ZN(n_0_0_68));
   AOI222_X1 i_0_0_106 (.A1(A[12]), .A2(n_0_0_119), .B1(n_0_0_96), .B2(A[16]), 
      .C1(A[20]), .C2(n_0_0_73), .ZN(n_0_0_69));
   OAI221_X1 i_0_0_107 (.A(n_0_0_70), .B1(n_0_0_101), .B2(n_0_0_75), .C1(
      n_0_0_71), .C2(n_0_0_100), .ZN(n_0_72));
   NAND2_X1 i_0_0_108 (.A1(A[13]), .A2(n_0_0_458), .ZN(n_0_0_70));
   MUX2_X1 i_0_0_109 (.A(n_0_0_80), .B(n_0_0_72), .S(n_0_0_125), .Z(n_0_0_71));
   AOI222_X1 i_0_0_110 (.A1(A[13]), .A2(n_0_0_119), .B1(n_0_0_96), .B2(A[17]), 
      .C1(A[21]), .C2(n_0_0_73), .ZN(n_0_0_72));
   AND2_X1 i_0_0_111 (.A1(n_0_0_84), .A2(n_0_0_462), .ZN(n_0_0_73));
   OAI221_X1 i_0_0_112 (.A(n_0_0_74), .B1(n_0_0_101), .B2(n_0_0_78), .C1(
      n_0_0_75), .C2(n_0_0_100), .ZN(n_0_73));
   NAND2_X1 i_0_0_113 (.A1(A[14]), .A2(n_0_0_458), .ZN(n_0_0_74));
   AOI222_X1 i_0_0_114 (.A1(n_0_0_76), .A2(n_0_0_125), .B1(A[16]), .B2(n_0_0_87), 
      .C1(n_0_0_97), .C2(n_0_0_96), .ZN(n_0_0_75));
   NOR2_X1 i_0_0_115 (.A1(n_0_0_77), .A2(n_0_0_124), .ZN(n_0_0_76));
   AOI22_X1 i_0_0_116 (.A1(A[14]), .A2(n_0_0_120), .B1(n_0_0_84), .B2(A[22]), 
      .ZN(n_0_0_77));
   OAI221_X1 i_0_0_117 (.A(n_0_0_85), .B1(n_0_0_78), .B2(n_0_0_100), .C1(
      n_0_0_86), .C2(n_0_0_101), .ZN(n_0_74));
   MUX2_X1 i_0_0_118 (.A(n_0_0_79), .B(n_0_0_80), .S(n_0_0_125), .Z(n_0_0_78));
   NAND2_X1 i_0_0_119 (.A1(n_0_0_120), .A2(n_0_0_92), .ZN(n_0_0_79));
   MUX2_X1 i_0_0_120 (.A(n_0_0_82), .B(n_0_0_81), .S(n_0_0_124), .Z(n_0_0_80));
   NAND2_X1 i_0_0_121 (.A1(A[19]), .A2(n_0_0_120), .ZN(n_0_0_81));
   OAI21_X1 i_0_0_122 (.A(n_0_0_123), .B1(n_0_0_121), .B2(A[15]), .ZN(n_0_0_82));
   NAND2_X1 i_0_0_123 (.A1(n_0_0_123), .A2(A[15]), .ZN(n_0_0_83));
   AND2_X1 i_0_0_124 (.A1(n_0_0_123), .A2(n_0_0_121), .ZN(n_0_0_84));
   NAND2_X1 i_0_0_125 (.A1(A[15]), .A2(n_0_0_458), .ZN(n_0_0_85));
   OAI221_X1 i_0_0_126 (.A(n_0_0_89), .B1(n_0_0_86), .B2(n_0_0_100), .C1(
      n_0_0_90), .C2(n_0_0_101), .ZN(n_0_75));
   AOI221_X1 i_0_0_127 (.A(n_0_0_88), .B1(n_0_0_87), .B2(A[18]), .C1(n_0_0_109), 
      .C2(n_0_0_96), .ZN(n_0_0_86));
   AND2_X1 i_0_0_128 (.A1(n_0_0_126), .A2(n_0_0_119), .ZN(n_0_0_87));
   AND3_X1 i_0_0_129 (.A1(A[16]), .A2(n_0_0_119), .A3(n_0_0_125), .ZN(n_0_0_88));
   NAND2_X1 i_0_0_130 (.A1(A[16]), .A2(n_0_0_458), .ZN(n_0_0_89));
   OAI221_X1 i_0_0_131 (.A(n_0_0_94), .B1(n_0_0_90), .B2(n_0_0_100), .C1(
      n_0_0_95), .C2(n_0_0_101), .ZN(n_0_76));
   OAI211_X1 i_0_0_132 (.A(n_0_0_120), .B(n_0_0_91), .C1(n_0_0_92), .C2(
      n_0_0_126), .ZN(n_0_0_90));
   OR3_X1 i_0_0_133 (.A1(n_0_0_125), .A2(n_0_0_124), .A3(A[19]), .ZN(n_0_0_91));
   OAI21_X1 i_0_0_134 (.A(n_0_0_93), .B1(n_0_0_462), .B2(n_0_0_441), .ZN(
      n_0_0_92));
   NAND2_X1 i_0_0_135 (.A1(n_0_0_462), .A2(A[17]), .ZN(n_0_0_93));
   NAND2_X1 i_0_0_136 (.A1(A[17]), .A2(n_0_0_458), .ZN(n_0_0_94));
   OAI221_X1 i_0_0_137 (.A(n_0_0_99), .B1(n_0_0_95), .B2(n_0_0_100), .C1(
      n_0_0_101), .C2(n_0_0_103), .ZN(n_0_77));
   AOI22_X1 i_0_0_138 (.A1(n_0_0_119), .A2(n_0_0_97), .B1(n_0_0_96), .B2(
      n_0_0_114), .ZN(n_0_0_95));
   NOR3_X1 i_0_0_139 (.A1(n_0_0_122), .A2(n_0_0_121), .A3(n_0_0_462), .ZN(
      n_0_0_96));
   OAI21_X1 i_0_0_140 (.A(n_0_0_98), .B1(n_0_0_125), .B2(n_0_0_440), .ZN(
      n_0_0_97));
   NAND2_X1 i_0_0_141 (.A1(n_0_0_125), .A2(A[18]), .ZN(n_0_0_98));
   NAND2_X1 i_0_0_142 (.A1(A[18]), .A2(n_0_0_458), .ZN(n_0_0_99));
   OAI221_X1 i_0_0_143 (.A(n_0_0_106), .B1(n_0_0_102), .B2(n_0_0_101), .C1(
      n_0_0_100), .C2(n_0_0_103), .ZN(n_0_78));
   NAND2_X1 i_0_0_144 (.A1(n_0_0_275), .A2(n_0_0_116), .ZN(n_0_0_100));
   NAND2_X1 i_0_0_145 (.A1(n_0_0_116), .A2(n_0_0_461), .ZN(n_0_0_101));
   NAND2_X1 i_0_0_146 (.A1(n_0_0_119), .A2(n_0_0_109), .ZN(n_0_0_102));
   AND2_X1 i_0_0_147 (.A1(n_0_0_105), .A2(n_0_0_104), .ZN(n_0_0_103));
   NAND3_X1 i_0_0_148 (.A1(A[21]), .A2(n_0_0_126), .A3(n_0_0_119), .ZN(n_0_0_104));
   OAI211_X1 i_0_0_149 (.A(n_0_0_120), .B(n_0_0_125), .C1(A[19]), .C2(n_0_0_124), 
      .ZN(n_0_0_105));
   NAND2_X1 i_0_0_150 (.A1(A[19]), .A2(n_0_0_458), .ZN(n_0_0_106));
   OAI22_X1 i_0_0_151 (.A1(n_0_0_115), .A2(n_0_0_107), .B1(n_0_0_440), .B2(
      n_0_0_410), .ZN(n_0_79));
   AOI21_X1 i_0_0_152 (.A(n_0_0_108), .B1(n_0_0_109), .B2(n_0_0_275), .ZN(
      n_0_0_107));
   NOR2_X1 i_0_0_153 (.A1(n_0_0_275), .A2(n_0_0_113), .ZN(n_0_0_108));
   OAI21_X1 i_0_0_154 (.A(n_0_0_110), .B1(n_0_0_126), .B2(n_0_0_440), .ZN(
      n_0_0_109));
   NAND2_X1 i_0_0_155 (.A1(A[22]), .A2(n_0_0_126), .ZN(n_0_0_110));
   OAI22_X1 i_0_0_156 (.A1(n_0_0_115), .A2(n_0_0_111), .B1(n_0_0_441), .B2(
      n_0_0_410), .ZN(n_0_80));
   AOI21_X1 i_0_0_157 (.A(n_0_0_112), .B1(n_0_0_114), .B2(n_0_0_461), .ZN(
      n_0_0_111));
   NOR2_X1 i_0_0_158 (.A1(n_0_0_113), .A2(n_0_0_461), .ZN(n_0_0_112));
   NOR2_X1 i_0_0_159 (.A1(A[21]), .A2(n_0_0_126), .ZN(n_0_0_113));
   AND2_X1 i_0_0_160 (.A1(n_0_0_125), .A2(A[22]), .ZN(n_0_0_114));
   NAND2_X1 i_0_0_161 (.A1(n_0_0_119), .A2(n_0_0_116), .ZN(n_0_0_115));
   AND2_X1 i_0_0_162 (.A1(n_0_0_410), .A2(n_0_0_127), .ZN(n_0_0_116));
   AOI21_X1 i_0_0_163 (.A(n_0_0_117), .B1(n_0_0_118), .B2(n_0_0_410), .ZN(n_0_81));
   AOI21_X1 i_0_0_164 (.A(A[22]), .B1(n_0_0_410), .B2(n_0_0_461), .ZN(n_0_0_117));
   NOR2_X1 i_0_0_165 (.A1(n_0_0_461), .A2(n_0_0_118), .ZN(n_0_82));
   NAND3_X1 i_0_0_166 (.A1(n_0_0_127), .A2(n_0_0_125), .A3(n_0_0_119), .ZN(
      n_0_0_118));
   NOR3_X1 i_0_0_167 (.A1(n_0_0_124), .A2(n_0_0_122), .A3(n_0_0_121), .ZN(
      n_0_0_119));
   NOR2_X1 i_0_0_168 (.A1(n_0_0_122), .A2(n_0_0_121), .ZN(n_0_0_120));
   XNOR2_X1 i_0_0_169 (.A(n_0_0_428), .B(n_0_0_257), .ZN(n_0_0_121));
   INV_X1 i_0_0_170 (.A(n_0_0_123), .ZN(n_0_0_122));
   XNOR2_X1 i_0_0_171 (.A(n_0_0_424), .B(n_0_0_260), .ZN(n_0_0_123));
   XOR2_X1 i_0_0_172 (.A(n_0_0_430), .B(n_0_0_254), .Z(n_0_0_124));
   XNOR2_X1 i_0_0_173 (.A(n_0_0_434), .B(n_0_0_250), .ZN(n_0_0_125));
   XNOR2_X1 i_0_0_174 (.A(n_0_0_433), .B(n_0_0_250), .ZN(n_0_0_126));
   AOI21_X1 i_0_0_175 (.A(n_0_0_128), .B1(n_0_0_263), .B2(n_0_0_419), .ZN(
      n_0_0_127));
   AOI221_X1 i_0_0_176 (.A(n_0_0_419), .B1(n_0_0_129), .B2(n_0_0_418), .C1(
      n_0_0_423), .C2(n_0_0_272), .ZN(n_0_0_128));
   MUX2_X1 i_0_0_177 (.A(n_0_0_414), .B(n_0_0_436), .S(n_0_0_273), .Z(n_0_0_129));
   OAI221_X1 i_0_0_178 (.A(n_0_0_133), .B1(n_0_0_130), .B2(n_0_0_244), .C1(
      n_0_0_224), .C2(n_0_0_134), .ZN(n_0_83));
   OAI21_X1 i_0_0_179 (.A(n_0_0_131), .B1(n_0_0_141), .B2(n_0_0_460), .ZN(
      n_0_0_130));
   OAI211_X1 i_0_0_180 (.A(n_0_0_132), .B(n_0_0_460), .C1(n_0_0_253), .C2(
      n_0_0_156), .ZN(n_0_0_131));
   AOI222_X1 i_0_0_181 (.A1(B[0]), .A2(n_0_0_252), .B1(n_0_0_207), .B2(B[8]), 
      .C1(B[16]), .C2(n_0_0_150), .ZN(n_0_0_132));
   NAND2_X1 i_0_0_182 (.A1(n_0_0_410), .A2(B[0]), .ZN(n_0_0_133));
   OAI221_X1 i_0_0_183 (.A(n_0_0_138), .B1(n_0_0_134), .B2(n_0_0_244), .C1(
      n_0_0_139), .C2(n_0_0_224), .ZN(n_0_84));
   OAI21_X1 i_0_0_184 (.A(n_0_0_137), .B1(n_0_0_135), .B2(n_0_0_249), .ZN(
      n_0_0_134));
   OAI21_X1 i_0_0_185 (.A(n_0_0_136), .B1(n_0_0_161), .B2(n_0_0_253), .ZN(
      n_0_0_135));
   AOI222_X1 i_0_0_186 (.A1(B[1]), .A2(n_0_0_252), .B1(n_0_0_207), .B2(B[9]), 
      .C1(B[17]), .C2(n_0_0_150), .ZN(n_0_0_136));
   NAND2_X1 i_0_0_187 (.A1(n_0_0_147), .A2(n_0_0_249), .ZN(n_0_0_137));
   NAND2_X1 i_0_0_188 (.A1(n_0_0_410), .A2(B[1]), .ZN(n_0_0_138));
   OAI221_X1 i_0_0_189 (.A(n_0_0_145), .B1(n_0_0_139), .B2(n_0_0_244), .C1(
      n_0_0_146), .C2(n_0_0_224), .ZN(n_0_85));
   OAI21_X1 i_0_0_190 (.A(n_0_0_140), .B1(n_0_0_141), .B2(n_0_0_249), .ZN(
      n_0_0_139));
   NAND2_X1 i_0_0_191 (.A1(n_0_0_154), .A2(n_0_0_249), .ZN(n_0_0_140));
   INV_X1 i_0_0_192 (.A(n_0_0_142), .ZN(n_0_0_141));
   AOI221_X1 i_0_0_193 (.A(n_0_0_143), .B1(n_0_0_168), .B2(n_0_0_459), .C1(B[18]), 
      .C2(n_0_0_150), .ZN(n_0_0_142));
   INV_X1 i_0_0_194 (.A(n_0_0_144), .ZN(n_0_0_143));
   AOI22_X1 i_0_0_195 (.A1(B[2]), .A2(n_0_0_252), .B1(n_0_0_207), .B2(B[10]), 
      .ZN(n_0_0_144));
   NAND2_X1 i_0_0_196 (.A1(n_0_0_410), .A2(B[2]), .ZN(n_0_0_145));
   OAI221_X1 i_0_0_197 (.A(n_0_0_151), .B1(n_0_0_224), .B2(n_0_0_152), .C1(
      n_0_0_146), .C2(n_0_0_244), .ZN(n_0_86));
   MUX2_X1 i_0_0_198 (.A(n_0_0_147), .B(n_0_0_159), .S(n_0_0_249), .Z(n_0_0_146));
   AOI221_X1 i_0_0_199 (.A(n_0_0_148), .B1(n_0_0_176), .B2(n_0_0_459), .C1(B[19]), 
      .C2(n_0_0_150), .ZN(n_0_0_147));
   INV_X1 i_0_0_200 (.A(n_0_0_149), .ZN(n_0_0_148));
   AOI22_X1 i_0_0_201 (.A1(B[3]), .A2(n_0_0_252), .B1(n_0_0_207), .B2(B[11]), 
      .ZN(n_0_0_149));
   NOR3_X1 i_0_0_202 (.A1(n_0_0_259), .A2(n_0_0_256), .A3(n_0_0_459), .ZN(
      n_0_0_150));
   NAND2_X1 i_0_0_203 (.A1(n_0_0_410), .A2(B[3]), .ZN(n_0_0_151));
   OAI221_X1 i_0_0_204 (.A(n_0_0_157), .B1(n_0_0_152), .B2(n_0_0_244), .C1(
      n_0_0_158), .C2(n_0_0_224), .ZN(n_0_87));
   OAI21_X1 i_0_0_205 (.A(n_0_0_153), .B1(n_0_0_165), .B2(n_0_0_460), .ZN(
      n_0_0_152));
   NAND2_X1 i_0_0_206 (.A1(n_0_0_460), .A2(n_0_0_154), .ZN(n_0_0_153));
   AOI221_X1 i_0_0_207 (.A(n_0_0_155), .B1(n_0_0_228), .B2(B[8]), .C1(B[16]), 
      .C2(n_0_0_187), .ZN(n_0_0_154));
   NOR2_X1 i_0_0_208 (.A1(n_0_0_459), .A2(n_0_0_156), .ZN(n_0_0_155));
   AOI222_X1 i_0_0_209 (.A1(B[4]), .A2(n_0_0_255), .B1(n_0_0_215), .B2(B[12]), 
      .C1(B[20]), .C2(n_0_0_171), .ZN(n_0_0_156));
   NAND2_X1 i_0_0_210 (.A1(n_0_0_410), .A2(B[4]), .ZN(n_0_0_157));
   OAI221_X1 i_0_0_211 (.A(n_0_0_162), .B1(n_0_0_224), .B2(n_0_0_163), .C1(
      n_0_0_158), .C2(n_0_0_244), .ZN(n_0_88));
   MUX2_X1 i_0_0_212 (.A(n_0_0_174), .B(n_0_0_159), .S(n_0_0_460), .Z(n_0_0_158));
   AOI221_X1 i_0_0_213 (.A(n_0_0_160), .B1(n_0_0_228), .B2(B[9]), .C1(B[17]), 
      .C2(n_0_0_187), .ZN(n_0_0_159));
   NOR2_X1 i_0_0_214 (.A1(n_0_0_459), .A2(n_0_0_161), .ZN(n_0_0_160));
   AOI222_X1 i_0_0_215 (.A1(B[5]), .A2(n_0_0_255), .B1(n_0_0_215), .B2(B[13]), 
      .C1(B[21]), .C2(n_0_0_171), .ZN(n_0_0_161));
   NAND2_X1 i_0_0_216 (.A1(n_0_0_410), .A2(B[5]), .ZN(n_0_0_162));
   OAI221_X1 i_0_0_217 (.A(n_0_0_172), .B1(n_0_0_163), .B2(n_0_0_244), .C1(
      n_0_0_224), .C2(n_0_0_173), .ZN(n_0_89));
   OAI21_X1 i_0_0_218 (.A(n_0_0_164), .B1(n_0_0_165), .B2(n_0_0_249), .ZN(
      n_0_0_163));
   NAND2_X1 i_0_0_219 (.A1(n_0_0_178), .A2(n_0_0_249), .ZN(n_0_0_164));
   NAND2_X1 i_0_0_220 (.A1(n_0_0_166), .A2(n_0_0_167), .ZN(n_0_0_165));
   AOI22_X1 i_0_0_221 (.A1(B[10]), .A2(n_0_0_228), .B1(n_0_0_187), .B2(B[18]), 
      .ZN(n_0_0_166));
   NAND2_X1 i_0_0_222 (.A1(n_0_0_253), .A2(n_0_0_168), .ZN(n_0_0_167));
   NAND2_X1 i_0_0_223 (.A1(n_0_0_169), .A2(n_0_0_170), .ZN(n_0_0_168));
   AOI22_X1 i_0_0_224 (.A1(B[14]), .A2(n_0_0_215), .B1(n_0_0_171), .B2(B[22]), 
      .ZN(n_0_0_169));
   NAND2_X1 i_0_0_225 (.A1(B[6]), .A2(n_0_0_255), .ZN(n_0_0_170));
   NOR2_X1 i_0_0_226 (.A1(n_0_0_259), .A2(n_0_0_256), .ZN(n_0_0_171));
   NAND2_X1 i_0_0_227 (.A1(n_0_0_410), .A2(B[6]), .ZN(n_0_0_172));
   OAI222_X1 i_0_0_228 (.A1(n_0_0_177), .A2(n_0_0_224), .B1(n_0_0_458), .B2(
      n_0_0_450), .C1(n_0_0_173), .C2(n_0_0_244), .ZN(n_0_90));
   MUX2_X1 i_0_0_229 (.A(n_0_0_181), .B(n_0_0_174), .S(n_0_0_460), .Z(n_0_0_173));
   AOI221_X1 i_0_0_230 (.A(n_0_0_175), .B1(n_0_0_176), .B2(n_0_0_253), .C1(B[19]), 
      .C2(n_0_0_187), .ZN(n_0_0_174));
   AND3_X1 i_0_0_231 (.A1(B[11]), .A2(n_0_0_255), .A3(n_0_0_459), .ZN(n_0_0_175));
   AOI22_X1 i_0_0_232 (.A1(n_0_0_255), .A2(n_0_0_450), .B1(n_0_0_256), .B2(
      n_0_0_214), .ZN(n_0_0_176));
   OAI221_X1 i_0_0_233 (.A(n_0_0_179), .B1(n_0_0_224), .B2(n_0_0_180), .C1(
      n_0_0_177), .C2(n_0_0_244), .ZN(n_0_91));
   MUX2_X1 i_0_0_234 (.A(n_0_0_184), .B(n_0_0_178), .S(n_0_0_460), .Z(n_0_0_177));
   AOI222_X1 i_0_0_235 (.A1(B[8]), .A2(n_0_0_252), .B1(n_0_0_196), .B2(n_0_0_459), 
      .C1(n_0_0_207), .C2(B[16]), .ZN(n_0_0_178));
   NAND2_X1 i_0_0_236 (.A1(n_0_0_410), .A2(B[8]), .ZN(n_0_0_179));
   OAI221_X1 i_0_0_237 (.A(n_0_0_182), .B1(n_0_0_180), .B2(n_0_0_244), .C1(
      n_0_0_224), .C2(n_0_0_183), .ZN(n_0_92));
   MUX2_X1 i_0_0_238 (.A(n_0_0_190), .B(n_0_0_181), .S(n_0_0_460), .Z(n_0_0_180));
   AOI222_X1 i_0_0_239 (.A1(B[9]), .A2(n_0_0_252), .B1(n_0_0_228), .B2(B[13]), 
      .C1(n_0_0_215), .C2(n_0_0_222), .ZN(n_0_0_181));
   NAND2_X1 i_0_0_240 (.A1(n_0_0_410), .A2(B[9]), .ZN(n_0_0_182));
   OAI221_X1 i_0_0_241 (.A(n_0_0_188), .B1(n_0_0_183), .B2(n_0_0_244), .C1(
      n_0_0_189), .C2(n_0_0_224), .ZN(n_0_93));
   MUX2_X1 i_0_0_242 (.A(n_0_0_195), .B(n_0_0_184), .S(n_0_0_460), .Z(n_0_0_183));
   AND2_X1 i_0_0_243 (.A1(n_0_0_186), .A2(n_0_0_185), .ZN(n_0_0_184));
   AOI22_X1 i_0_0_244 (.A1(B[10]), .A2(n_0_0_252), .B1(n_0_0_228), .B2(B[14]), 
      .ZN(n_0_0_185));
   AOI22_X1 i_0_0_245 (.A1(B[18]), .A2(n_0_0_207), .B1(n_0_0_187), .B2(B[22]), 
      .ZN(n_0_0_186));
   AND2_X1 i_0_0_246 (.A1(n_0_0_459), .A2(n_0_0_215), .ZN(n_0_0_187));
   NAND2_X1 i_0_0_247 (.A1(n_0_0_410), .A2(B[10]), .ZN(n_0_0_188));
   OAI221_X1 i_0_0_248 (.A(n_0_0_193), .B1(n_0_0_189), .B2(n_0_0_244), .C1(
      n_0_0_224), .C2(n_0_0_194), .ZN(n_0_94));
   MUX2_X1 i_0_0_249 (.A(n_0_0_190), .B(n_0_0_201), .S(n_0_0_249), .Z(n_0_0_189));
   OAI211_X1 i_0_0_250 (.A(n_0_0_259), .B(n_0_0_192), .C1(n_0_0_191), .C2(
      n_0_0_256), .ZN(n_0_0_190));
   MUX2_X1 i_0_0_251 (.A(B[11]), .B(B[15]), .S(n_0_0_459), .Z(n_0_0_191));
   NAND2_X1 i_0_0_252 (.A1(n_0_0_256), .A2(n_0_0_236), .ZN(n_0_0_192));
   NAND2_X1 i_0_0_253 (.A1(n_0_0_410), .A2(B[11]), .ZN(n_0_0_193));
   OAI221_X1 i_0_0_254 (.A(n_0_0_198), .B1(n_0_0_224), .B2(n_0_0_199), .C1(
      n_0_0_194), .C2(n_0_0_244), .ZN(n_0_95));
   MUX2_X1 i_0_0_255 (.A(n_0_0_195), .B(n_0_0_206), .S(n_0_0_249), .Z(n_0_0_194));
   AOI22_X1 i_0_0_256 (.A1(n_0_0_196), .A2(n_0_0_253), .B1(B[16]), .B2(n_0_0_228), 
      .ZN(n_0_0_195));
   INV_X1 i_0_0_257 (.A(n_0_0_197), .ZN(n_0_0_196));
   AOI22_X1 i_0_0_258 (.A1(B[12]), .A2(n_0_0_255), .B1(n_0_0_215), .B2(B[20]), 
      .ZN(n_0_0_197));
   NAND2_X1 i_0_0_259 (.A1(n_0_0_410), .A2(B[12]), .ZN(n_0_0_198));
   OAI221_X1 i_0_0_260 (.A(n_0_0_202), .B1(n_0_0_199), .B2(n_0_0_244), .C1(
      n_0_0_203), .C2(n_0_0_224), .ZN(n_0_96));
   OAI21_X1 i_0_0_261 (.A(n_0_0_200), .B1(n_0_0_211), .B2(n_0_0_460), .ZN(
      n_0_0_199));
   NAND2_X1 i_0_0_262 (.A1(n_0_0_460), .A2(n_0_0_201), .ZN(n_0_0_200));
   AOI222_X1 i_0_0_263 (.A1(B[13]), .A2(n_0_0_252), .B1(n_0_0_228), .B2(B[17]), 
      .C1(B[21]), .C2(n_0_0_207), .ZN(n_0_0_201));
   NAND2_X1 i_0_0_264 (.A1(n_0_0_410), .A2(B[13]), .ZN(n_0_0_202));
   OAI221_X1 i_0_0_265 (.A(n_0_0_208), .B1(n_0_0_224), .B2(n_0_0_209), .C1(
      n_0_0_203), .C2(n_0_0_244), .ZN(n_0_97));
   AOI21_X1 i_0_0_266 (.A(n_0_0_204), .B1(n_0_0_226), .B2(B[16]), .ZN(n_0_0_203));
   OAI21_X1 i_0_0_267 (.A(n_0_0_205), .B1(n_0_0_206), .B2(n_0_0_249), .ZN(
      n_0_0_204));
   NAND3_X1 i_0_0_268 (.A1(B[20]), .A2(n_0_0_249), .A3(n_0_0_228), .ZN(n_0_0_205));
   AOI222_X1 i_0_0_269 (.A1(B[14]), .A2(n_0_0_252), .B1(n_0_0_228), .B2(B[18]), 
      .C1(B[22]), .C2(n_0_0_207), .ZN(n_0_0_206));
   AND2_X1 i_0_0_270 (.A1(n_0_0_215), .A2(n_0_0_253), .ZN(n_0_0_207));
   NAND2_X1 i_0_0_271 (.A1(n_0_0_410), .A2(B[14]), .ZN(n_0_0_208));
   OAI221_X1 i_0_0_272 (.A(n_0_0_216), .B1(n_0_0_244), .B2(n_0_0_209), .C1(
      n_0_0_217), .C2(n_0_0_224), .ZN(n_0_98));
   AOI21_X1 i_0_0_273 (.A(n_0_0_210), .B1(n_0_0_211), .B2(n_0_0_460), .ZN(
      n_0_0_209));
   AND3_X1 i_0_0_274 (.A1(n_0_0_255), .A2(n_0_0_249), .A3(n_0_0_222), .ZN(
      n_0_0_210));
   OAI21_X1 i_0_0_275 (.A(n_0_0_212), .B1(n_0_0_213), .B2(n_0_0_459), .ZN(
      n_0_0_211));
   NAND3_X1 i_0_0_276 (.A1(B[19]), .A2(n_0_0_255), .A3(n_0_0_459), .ZN(n_0_0_212));
   OAI21_X1 i_0_0_277 (.A(n_0_0_259), .B1(n_0_0_256), .B2(B[15]), .ZN(n_0_0_213));
   NAND2_X1 i_0_0_278 (.A1(n_0_0_259), .A2(B[15]), .ZN(n_0_0_214));
   AND2_X1 i_0_0_279 (.A1(n_0_0_259), .A2(n_0_0_256), .ZN(n_0_0_215));
   NAND2_X1 i_0_0_280 (.A1(n_0_0_410), .A2(B[15]), .ZN(n_0_0_216));
   OAI221_X1 i_0_0_281 (.A(n_0_0_219), .B1(n_0_0_217), .B2(n_0_0_244), .C1(
      n_0_0_224), .C2(n_0_0_220), .ZN(n_0_99));
   AOI221_X1 i_0_0_282 (.A(n_0_0_218), .B1(n_0_0_248), .B2(B[16]), .C1(B[18]), 
      .C2(n_0_0_226), .ZN(n_0_0_217));
   AND2_X1 i_0_0_283 (.A1(n_0_0_228), .A2(n_0_0_240), .ZN(n_0_0_218));
   NAND2_X1 i_0_0_284 (.A1(n_0_0_410), .A2(B[16]), .ZN(n_0_0_219));
   OAI221_X1 i_0_0_285 (.A(n_0_0_223), .B1(n_0_0_220), .B2(n_0_0_244), .C1(
      n_0_0_225), .C2(n_0_0_224), .ZN(n_0_100));
   OAI211_X1 i_0_0_286 (.A(n_0_0_255), .B(n_0_0_221), .C1(n_0_0_222), .C2(
      n_0_0_249), .ZN(n_0_0_220));
   NAND2_X1 i_0_0_287 (.A1(n_0_0_249), .A2(n_0_0_236), .ZN(n_0_0_221));
   MUX2_X1 i_0_0_288 (.A(B[17]), .B(B[21]), .S(n_0_0_459), .Z(n_0_0_222));
   NAND2_X1 i_0_0_289 (.A1(n_0_0_410), .A2(B[17]), .ZN(n_0_0_223));
   OAI221_X1 i_0_0_290 (.A(n_0_0_229), .B1(n_0_0_225), .B2(n_0_0_244), .C1(
      n_0_0_224), .C2(n_0_0_233), .ZN(n_0_101));
   NAND2_X1 i_0_0_291 (.A1(n_0_0_245), .A2(n_0_0_461), .ZN(n_0_0_224));
   AOI221_X1 i_0_0_292 (.A(n_0_0_227), .B1(n_0_0_226), .B2(B[20]), .C1(B[18]), 
      .C2(n_0_0_248), .ZN(n_0_0_225));
   NOR2_X1 i_0_0_293 (.A1(n_0_0_251), .A2(n_0_0_460), .ZN(n_0_0_226));
   AND3_X1 i_0_0_294 (.A1(B[22]), .A2(n_0_0_228), .A3(n_0_0_460), .ZN(n_0_0_227));
   NOR3_X1 i_0_0_295 (.A1(n_0_0_258), .A2(n_0_0_256), .A3(n_0_0_253), .ZN(
      n_0_0_228));
   NAND2_X1 i_0_0_296 (.A1(n_0_0_410), .A2(B[18]), .ZN(n_0_0_229));
   INV_X1 i_0_0_297 (.A(n_0_0_230), .ZN(n_0_102));
   AOI22_X1 i_0_0_298 (.A1(n_0_0_231), .A2(n_0_0_245), .B1(n_0_0_410), .B2(B[19]), 
      .ZN(n_0_0_230));
   OAI21_X1 i_0_0_299 (.A(n_0_0_232), .B1(n_0_0_233), .B2(n_0_0_461), .ZN(
      n_0_0_231));
   NAND3_X1 i_0_0_300 (.A1(n_0_0_252), .A2(n_0_0_240), .A3(n_0_0_461), .ZN(
      n_0_0_232));
   NAND2_X1 i_0_0_301 (.A1(n_0_0_255), .A2(n_0_0_234), .ZN(n_0_0_233));
   OAI21_X1 i_0_0_302 (.A(n_0_0_235), .B1(n_0_0_236), .B2(n_0_0_249), .ZN(
      n_0_0_234));
   NAND3_X1 i_0_0_303 (.A1(n_0_0_253), .A2(n_0_0_249), .A3(B[21]), .ZN(n_0_0_235));
   NOR2_X1 i_0_0_304 (.A1(B[19]), .A2(n_0_0_459), .ZN(n_0_0_236));
   OAI21_X1 i_0_0_305 (.A(n_0_0_237), .B1(n_0_0_458), .B2(n_0_0_451), .ZN(
      n_0_103));
   NAND3_X1 i_0_0_306 (.A1(n_0_0_252), .A2(n_0_0_245), .A3(n_0_0_238), .ZN(
      n_0_0_237));
   AOI21_X1 i_0_0_307 (.A(n_0_0_239), .B1(n_0_0_241), .B2(n_0_0_275), .ZN(
      n_0_0_238));
   NOR3_X1 i_0_0_308 (.A1(B[21]), .A2(n_0_0_275), .A3(n_0_0_249), .ZN(n_0_0_239));
   INV_X1 i_0_0_309 (.A(n_0_0_241), .ZN(n_0_0_240));
   AOI21_X1 i_0_0_310 (.A(n_0_0_242), .B1(n_0_0_249), .B2(B[22]), .ZN(n_0_0_241));
   NOR2_X1 i_0_0_311 (.A1(n_0_0_249), .A2(n_0_0_451), .ZN(n_0_0_242));
   OAI211_X1 i_0_0_312 (.A(n_0_0_246), .B(n_0_0_243), .C1(n_0_0_244), .C2(
      n_0_0_251), .ZN(n_0_104));
   NAND3_X1 i_0_0_313 (.A1(B[22]), .A2(n_0_0_248), .A3(n_0_0_245), .ZN(n_0_0_243));
   NAND2_X1 i_0_0_314 (.A1(n_0_0_275), .A2(n_0_0_245), .ZN(n_0_0_244));
   NOR2_X1 i_0_0_315 (.A1(n_0_0_410), .A2(n_0_0_262), .ZN(n_0_0_245));
   NAND2_X1 i_0_0_316 (.A1(n_0_0_410), .A2(B[21]), .ZN(n_0_0_246));
   NOR2_X1 i_0_0_317 (.A1(n_0_0_274), .A2(n_0_0_247), .ZN(n_0_105));
   AOI21_X1 i_0_0_318 (.A(n_0_0_410), .B1(n_0_0_261), .B2(n_0_0_248), .ZN(
      n_0_0_247));
   NOR2_X1 i_0_0_319 (.A1(n_0_0_251), .A2(n_0_0_249), .ZN(n_0_0_248));
   XOR2_X1 i_0_0_320 (.A(n_0_0_276), .B(n_0_0_250), .Z(n_0_0_249));
   XNOR2_X1 i_0_0_321 (.A(n_0_0_453), .B(A[24]), .ZN(n_0_0_250));
   NAND2_X1 i_0_0_322 (.A1(n_0_0_255), .A2(n_0_0_253), .ZN(n_0_0_251));
   NOR3_X1 i_0_0_323 (.A1(n_0_0_258), .A2(n_0_0_256), .A3(n_0_0_459), .ZN(
      n_0_0_252));
   XOR2_X1 i_0_0_324 (.A(n_0_0_269), .B(n_0_0_254), .Z(n_0_0_253));
   XNOR2_X1 i_0_0_325 (.A(B[25]), .B(n_0_0_443), .ZN(n_0_0_254));
   NOR2_X1 i_0_0_326 (.A1(n_0_0_258), .A2(n_0_0_256), .ZN(n_0_0_255));
   XOR2_X1 i_0_0_327 (.A(n_0_0_268), .B(n_0_0_257), .Z(n_0_0_256));
   NAND2_X1 i_0_0_328 (.A1(n_0_0_426), .A2(n_0_0_425), .ZN(n_0_0_257));
   INV_X1 i_0_0_329 (.A(n_0_0_259), .ZN(n_0_0_258));
   XNOR2_X1 i_0_0_330 (.A(n_0_0_266), .B(n_0_0_260), .ZN(n_0_0_259));
   XNOR2_X1 i_0_0_331 (.A(B[27]), .B(n_0_0_445), .ZN(n_0_0_260));
   INV_X1 i_0_0_332 (.A(n_0_0_262), .ZN(n_0_0_261));
   MUX2_X1 i_0_0_333 (.A(n_0_0_263), .B(n_0_0_270), .S(n_0_0_264), .Z(n_0_0_262));
   NAND3_X1 i_0_0_334 (.A1(n_0_0_272), .A2(n_0_0_417), .A3(n_0_0_422), .ZN(
      n_0_0_263));
   AOI21_X1 i_0_0_335 (.A(n_0_0_420), .B1(n_0_0_265), .B2(n_0_0_421), .ZN(
      n_0_0_264));
   INV_X1 i_0_0_336 (.A(n_0_0_266), .ZN(n_0_0_265));
   AOI21_X1 i_0_0_337 (.A(n_0_0_267), .B1(A[26]), .B2(n_0_0_454), .ZN(n_0_0_266));
   NOR2_X1 i_0_0_338 (.A1(n_0_0_427), .A2(n_0_0_268), .ZN(n_0_0_267));
   OAI21_X1 i_0_0_339 (.A(n_0_0_429), .B1(n_0_0_269), .B2(n_0_0_435), .ZN(
      n_0_0_268));
   OAI21_X1 i_0_0_340 (.A(n_0_0_431), .B1(n_0_0_276), .B2(n_0_0_432), .ZN(
      n_0_0_269));
   AOI22_X1 i_0_0_341 (.A1(n_0_0_271), .A2(n_0_0_423), .B1(n_0_0_418), .B2(
      n_0_0_272), .ZN(n_0_0_270));
   MUX2_X1 i_0_0_342 (.A(n_0_0_436), .B(n_0_0_414), .S(n_0_0_273), .Z(n_0_0_271));
   NOR3_X1 i_0_0_343 (.A1(n_0_0_273), .A2(n_0_0_414), .A3(n_0_0_436), .ZN(
      n_0_0_272));
   NAND2_X1 i_0_0_344 (.A1(n_0_0_413), .A2(n_0_0_412), .ZN(n_0_0_273));
   AOI21_X1 i_0_0_345 (.A(B[22]), .B1(n_0_0_458), .B2(n_0_0_461), .ZN(n_0_0_274));
   NOR2_X1 i_0_0_346 (.A1(n_0_0_434), .A2(n_0_0_276), .ZN(n_0_0_275));
   NOR2_X1 i_0_0_347 (.A1(n_0_0_452), .A2(A[23]), .ZN(n_0_0_276));
   AND2_X1 i_0_0_348 (.A1(n_0_25), .A2(n_0_111), .ZN(n_0_107));
   AND2_X1 i_0_0_349 (.A1(n_0_26), .A2(n_0_111), .ZN(n_0_108));
   AND2_X1 i_0_0_350 (.A1(n_0_27), .A2(n_0_111), .ZN(n_0_109));
   AND2_X1 i_0_0_351 (.A1(n_0_28), .A2(n_0_111), .ZN(n_0_110));
   AND2_X1 i_0_0_352 (.A1(n_0_29), .A2(n_0_111), .ZN(n_0_112));
   NOR3_X1 i_0_0_353 (.A1(n_0_0_278), .A2(n_0_0_277), .A3(A[31]), .ZN(overflow));
   NOR3_X1 i_0_0_354 (.A1(n_0_0_449), .A2(n_0_0_278), .A3(n_0_0_277), .ZN(
      underflow));
   OAI211_X1 i_0_0_355 (.A(n_0_114), .B(n_0_0_282), .C1(n_0_0_442), .C2(
      n_0_0_410), .ZN(n_0_0_277));
   NAND4_X1 i_0_0_356 (.A1(n_0_0_279), .A2(n_0_115), .A3(n_0_116), .A4(n_0_117), 
      .ZN(n_0_0_278));
   AOI221_X1 i_0_0_357 (.A(n_0_0_403), .B1(n_0_0_281), .B2(n_0_0_280), .C1(
      n_0_0_448), .C2(n_0_0_456), .ZN(n_0_0_279));
   NAND3_X1 i_0_0_358 (.A1(n_0_0_410), .A2(B[28]), .A3(B[29]), .ZN(n_0_0_280));
   NAND3_X1 i_0_0_359 (.A1(A[29]), .A2(A[28]), .A3(n_0_0_458), .ZN(n_0_0_281));
   OAI21_X1 i_0_0_360 (.A(n_0_0_282), .B1(n_0_0_410), .B2(n_0_0_442), .ZN(
      n_0_113));
   NAND2_X1 i_0_0_361 (.A1(n_0_0_410), .A2(B[23]), .ZN(n_0_0_282));
   OAI21_X1 i_0_0_362 (.A(n_0_0_283), .B1(n_0_0_458), .B2(n_0_0_453), .ZN(
      n_0_114));
   NAND2_X1 i_0_0_363 (.A1(A[24]), .A2(n_0_0_458), .ZN(n_0_0_283));
   OAI21_X1 i_0_0_364 (.A(n_0_0_284), .B1(n_0_0_410), .B2(n_0_0_443), .ZN(
      n_0_115));
   NAND2_X1 i_0_0_365 (.A1(n_0_0_410), .A2(B[25]), .ZN(n_0_0_284));
   OAI21_X1 i_0_0_366 (.A(n_0_0_285), .B1(n_0_0_410), .B2(n_0_0_444), .ZN(
      n_0_116));
   NAND2_X1 i_0_0_367 (.A1(n_0_0_410), .A2(B[26]), .ZN(n_0_0_285));
   OAI21_X1 i_0_0_368 (.A(n_0_0_286), .B1(n_0_0_410), .B2(n_0_0_445), .ZN(
      n_0_117));
   NAND2_X1 i_0_0_369 (.A1(n_0_0_410), .A2(B[27]), .ZN(n_0_0_286));
   OAI21_X1 i_0_0_370 (.A(n_0_0_287), .B1(n_0_0_410), .B2(n_0_0_446), .ZN(
      n_0_118));
   NAND2_X1 i_0_0_371 (.A1(n_0_0_410), .A2(B[28]), .ZN(n_0_0_287));
   OAI21_X1 i_0_0_372 (.A(n_0_0_288), .B1(n_0_0_410), .B2(n_0_0_447), .ZN(
      n_0_119));
   NAND2_X1 i_0_0_373 (.A1(n_0_0_410), .A2(B[29]), .ZN(n_0_0_288));
   NAND2_X1 i_0_0_374 (.A1(n_0_0_456), .A2(n_0_0_448), .ZN(n_0_120));
   NOR2_X1 i_0_0_375 (.A1(n_0_0_290), .A2(n_0_0_289), .ZN(Sum[0]));
   AOI21_X1 i_0_0_376 (.A(n_0_0_404), .B1(n_0_0_305), .B2(num_leading_zeros[0]), 
      .ZN(n_0_0_289));
   INV_X1 i_0_0_377 (.A(n_0_0_291), .ZN(n_0_0_290));
   OAI21_X1 i_0_0_378 (.A(n_0_0_292), .B1(n_0_0_403), .B2(n_0_0_438), .ZN(
      n_0_0_291));
   NAND2_X1 i_0_0_379 (.A1(n_0_0_403), .A2(n_0_0), .ZN(n_0_0_292));
   AOI21_X1 i_0_0_380 (.A(n_0_0_293), .B1(n_0_0_296), .B2(n_0_0_408), .ZN(Sum[1]));
   AOI221_X1 i_0_0_381 (.A(n_0_0_408), .B1(n_0_0_405), .B2(n_0_1), .C1(n_0_0_305), 
      .C2(n_0_0_294), .ZN(n_0_0_293));
   OAI21_X1 i_0_0_382 (.A(n_0_0_295), .B1(n_0_0_438), .B2(n_0_57), .ZN(n_0_0_294));
   NAND3_X1 i_0_0_383 (.A1(n_0_57), .A2(n_0_0_406), .A3(n_0_0), .ZN(n_0_0_295));
   AOI21_X1 i_0_0_384 (.A(n_0_0_297), .B1(n_0_2), .B2(n_0_24), .ZN(n_0_0_296));
   NOR2_X1 i_0_0_385 (.A1(n_0_0_438), .A2(n_0_24), .ZN(n_0_0_297));
   NOR2_X1 i_0_0_386 (.A1(n_0_0_299), .A2(n_0_0_298), .ZN(Sum[2]));
   OAI22_X1 i_0_0_387 (.A1(n_0_106), .A2(n_0_2), .B1(n_0_3), .B2(n_0_0_403), 
      .ZN(n_0_0_298));
   NOR2_X1 i_0_0_388 (.A1(n_0_0_300), .A2(n_0_0_404), .ZN(n_0_0_299));
   AOI21_X1 i_0_0_389 (.A(n_0_0_301), .B1(n_0_0_302), .B2(num_leading_zeros[0]), 
      .ZN(n_0_0_300));
   AOI21_X1 i_0_0_390 (.A(num_leading_zeros[0]), .B1(n_0_1), .B2(n_0_0_305), 
      .ZN(n_0_0_301));
   AOI221_X1 i_0_0_391 (.A(n_0_0_303), .B1(n_0_0_302), .B2(n_0_0_363), .C1(
      n_0_0_304), .C2(n_0_0_364), .ZN(Sum[3]));
   AOI22_X1 i_0_0_392 (.A1(n_0_0), .A2(n_0_0_312), .B1(n_0_0_305), .B2(n_0_2), 
      .ZN(n_0_0_302));
   OAI22_X1 i_0_0_393 (.A1(n_0_106), .A2(n_0_3), .B1(n_0_4), .B2(n_0_0_403), 
      .ZN(n_0_0_303));
   AOI221_X1 i_0_0_394 (.A(n_0_0_306), .B1(n_0_0_304), .B2(n_0_0_363), .C1(
      n_0_0_307), .C2(n_0_0_364), .ZN(Sum[4]));
   AOI22_X1 i_0_0_395 (.A1(n_0_1), .A2(n_0_0_312), .B1(n_0_0_305), .B2(n_0_3), 
      .ZN(n_0_0_304));
   NOR3_X1 i_0_0_396 (.A1(n_0_0_398), .A2(n_0_58), .A3(n_0_59), .ZN(n_0_0_305));
   OAI22_X1 i_0_0_397 (.A1(n_0_106), .A2(n_0_4), .B1(n_0_5), .B2(n_0_0_403), 
      .ZN(n_0_0_306));
   AOI221_X1 i_0_0_398 (.A(n_0_0_309), .B1(n_0_0_307), .B2(n_0_0_363), .C1(
      n_0_0_310), .C2(n_0_0_364), .ZN(Sum[5]));
   AOI21_X1 i_0_0_399 (.A(n_0_0_308), .B1(n_0_0_312), .B2(n_0_2), .ZN(n_0_0_307));
   NOR2_X1 i_0_0_400 (.A1(n_0_0_315), .A2(n_0_58), .ZN(n_0_0_308));
   OAI22_X1 i_0_0_401 (.A1(n_0_106), .A2(n_0_5), .B1(n_0_6), .B2(n_0_0_403), 
      .ZN(n_0_0_309));
   AOI221_X1 i_0_0_402 (.A(n_0_0_313), .B1(n_0_0_310), .B2(n_0_0_363), .C1(
      n_0_0_314), .C2(n_0_0_364), .ZN(Sum[6]));
   AOI21_X1 i_0_0_403 (.A(n_0_0_311), .B1(n_0_0_312), .B2(n_0_3), .ZN(n_0_0_310));
   NOR2_X1 i_0_0_404 (.A1(n_0_0_318), .A2(n_0_58), .ZN(n_0_0_311));
   AND2_X1 i_0_0_405 (.A1(n_0_58), .A2(n_0_0_394), .ZN(n_0_0_312));
   OAI22_X1 i_0_0_406 (.A1(n_0_106), .A2(n_0_6), .B1(n_0_7), .B2(n_0_0_403), 
      .ZN(n_0_0_313));
   AOI221_X1 i_0_0_407 (.A(n_0_0_316), .B1(n_0_0_314), .B2(n_0_0_363), .C1(
      n_0_0_317), .C2(n_0_0_364), .ZN(Sum[7]));
   MUX2_X1 i_0_0_408 (.A(n_0_0_321), .B(n_0_0_315), .S(n_0_58), .Z(n_0_0_314));
   AOI22_X1 i_0_0_409 (.A1(n_0_4), .A2(n_0_0_394), .B1(n_0_0_353), .B2(n_0_0), 
      .ZN(n_0_0_315));
   OAI22_X1 i_0_0_410 (.A1(n_0_106), .A2(n_0_7), .B1(n_0_8), .B2(n_0_0_403), 
      .ZN(n_0_0_316));
   AOI221_X1 i_0_0_411 (.A(n_0_0_319), .B1(n_0_0_317), .B2(n_0_0_363), .C1(
      n_0_0_320), .C2(n_0_0_364), .ZN(Sum[8]));
   MUX2_X1 i_0_0_412 (.A(n_0_0_324), .B(n_0_0_318), .S(n_0_58), .Z(n_0_0_317));
   AOI22_X1 i_0_0_413 (.A1(n_0_5), .A2(n_0_0_394), .B1(n_0_0_353), .B2(n_0_1), 
      .ZN(n_0_0_318));
   OAI22_X1 i_0_0_414 (.A1(n_0_106), .A2(n_0_8), .B1(n_0_9), .B2(n_0_0_403), 
      .ZN(n_0_0_319));
   AOI221_X1 i_0_0_415 (.A(n_0_0_322), .B1(n_0_0_320), .B2(n_0_0_363), .C1(
      n_0_0_323), .C2(n_0_0_364), .ZN(Sum[9]));
   MUX2_X1 i_0_0_416 (.A(n_0_0_327), .B(n_0_0_321), .S(n_0_58), .Z(n_0_0_320));
   AOI22_X1 i_0_0_417 (.A1(n_0_6), .A2(n_0_0_394), .B1(n_0_0_353), .B2(n_0_2), 
      .ZN(n_0_0_321));
   OAI22_X1 i_0_0_418 (.A1(n_0_106), .A2(n_0_9), .B1(n_0_10), .B2(n_0_0_403), 
      .ZN(n_0_0_322));
   AOI221_X1 i_0_0_419 (.A(n_0_0_325), .B1(n_0_0_323), .B2(n_0_0_363), .C1(
      n_0_0_326), .C2(n_0_0_364), .ZN(Sum[10]));
   MUX2_X1 i_0_0_420 (.A(n_0_0_330), .B(n_0_0_324), .S(n_0_58), .Z(n_0_0_323));
   AOI22_X1 i_0_0_421 (.A1(n_0_7), .A2(n_0_0_394), .B1(n_0_0_353), .B2(n_0_3), 
      .ZN(n_0_0_324));
   OAI22_X1 i_0_0_422 (.A1(n_0_106), .A2(n_0_10), .B1(n_0_11), .B2(n_0_0_403), 
      .ZN(n_0_0_325));
   AOI221_X1 i_0_0_423 (.A(n_0_0_328), .B1(n_0_0_326), .B2(n_0_0_363), .C1(
      n_0_0_329), .C2(n_0_0_364), .ZN(Sum[11]));
   MUX2_X1 i_0_0_424 (.A(n_0_0_333), .B(n_0_0_327), .S(n_0_58), .Z(n_0_0_326));
   AOI222_X1 i_0_0_425 (.A1(n_0_8), .A2(n_0_0_394), .B1(n_0_0_392), .B2(n_0_0), 
      .C1(n_0_0_353), .C2(n_0_4), .ZN(n_0_0_327));
   OAI22_X1 i_0_0_426 (.A1(n_0_106), .A2(n_0_11), .B1(n_0_12), .B2(n_0_0_403), 
      .ZN(n_0_0_328));
   AOI221_X1 i_0_0_427 (.A(n_0_0_331), .B1(n_0_0_329), .B2(n_0_0_363), .C1(
      n_0_0_332), .C2(n_0_0_364), .ZN(Sum[12]));
   MUX2_X1 i_0_0_428 (.A(n_0_0_336), .B(n_0_0_330), .S(n_0_58), .Z(n_0_0_329));
   AOI222_X1 i_0_0_429 (.A1(n_0_9), .A2(n_0_0_394), .B1(n_0_0_392), .B2(n_0_1), 
      .C1(n_0_0_353), .C2(n_0_5), .ZN(n_0_0_330));
   OAI22_X1 i_0_0_430 (.A1(n_0_106), .A2(n_0_12), .B1(n_0_13), .B2(n_0_0_403), 
      .ZN(n_0_0_331));
   AOI221_X1 i_0_0_431 (.A(n_0_0_334), .B1(n_0_0_332), .B2(n_0_0_363), .C1(
      n_0_0_335), .C2(n_0_0_364), .ZN(Sum[13]));
   MUX2_X1 i_0_0_432 (.A(n_0_0_339), .B(n_0_0_333), .S(n_0_58), .Z(n_0_0_332));
   AOI222_X1 i_0_0_433 (.A1(n_0_10), .A2(n_0_0_394), .B1(n_0_0_392), .B2(n_0_2), 
      .C1(n_0_0_353), .C2(n_0_6), .ZN(n_0_0_333));
   OAI22_X1 i_0_0_434 (.A1(n_0_106), .A2(n_0_13), .B1(n_0_14), .B2(n_0_0_403), 
      .ZN(n_0_0_334));
   AOI221_X1 i_0_0_435 (.A(n_0_0_337), .B1(n_0_0_335), .B2(n_0_0_363), .C1(
      n_0_0_338), .C2(n_0_0_364), .ZN(Sum[14]));
   MUX2_X1 i_0_0_436 (.A(n_0_0_343), .B(n_0_0_336), .S(n_0_58), .Z(n_0_0_335));
   AOI222_X1 i_0_0_437 (.A1(n_0_11), .A2(n_0_0_394), .B1(n_0_0_392), .B2(n_0_3), 
      .C1(n_0_0_353), .C2(n_0_7), .ZN(n_0_0_336));
   OAI22_X1 i_0_0_438 (.A1(n_0_106), .A2(n_0_14), .B1(n_0_15), .B2(n_0_0_403), 
      .ZN(n_0_0_337));
   AOI221_X1 i_0_0_439 (.A(n_0_0_341), .B1(n_0_0_338), .B2(n_0_0_363), .C1(
      n_0_0_342), .C2(n_0_0_364), .ZN(Sum[15]));
   MUX2_X1 i_0_0_440 (.A(n_0_0_347), .B(n_0_0_339), .S(n_0_58), .Z(n_0_0_338));
   AOI221_X1 i_0_0_441 (.A(n_0_0_340), .B1(n_0_0_352), .B2(n_0_0), .C1(n_0_8), 
      .C2(n_0_0_353), .ZN(n_0_0_339));
   NOR2_X1 i_0_0_442 (.A1(n_0_0_357), .A2(n_0_59), .ZN(n_0_0_340));
   OAI22_X1 i_0_0_443 (.A1(n_0_106), .A2(n_0_15), .B1(n_0_16), .B2(n_0_0_403), 
      .ZN(n_0_0_341));
   AOI221_X1 i_0_0_444 (.A(n_0_0_345), .B1(n_0_0_342), .B2(n_0_0_363), .C1(
      n_0_0_346), .C2(n_0_0_364), .ZN(Sum[16]));
   MUX2_X1 i_0_0_445 (.A(n_0_0_351), .B(n_0_0_343), .S(n_0_58), .Z(n_0_0_342));
   AOI221_X1 i_0_0_446 (.A(n_0_0_344), .B1(n_0_0_352), .B2(n_0_1), .C1(n_0_9), 
      .C2(n_0_0_353), .ZN(n_0_0_343));
   NOR2_X1 i_0_0_447 (.A1(n_0_0_361), .A2(n_0_59), .ZN(n_0_0_344));
   OAI22_X1 i_0_0_448 (.A1(n_0_106), .A2(n_0_16), .B1(n_0_17), .B2(n_0_0_403), 
      .ZN(n_0_0_345));
   AOI221_X1 i_0_0_449 (.A(n_0_0_349), .B1(n_0_0_364), .B2(n_0_0_350), .C1(
      n_0_0_346), .C2(n_0_0_363), .ZN(Sum[17]));
   MUX2_X1 i_0_0_450 (.A(n_0_0_356), .B(n_0_0_347), .S(n_0_58), .Z(n_0_0_346));
   AOI221_X1 i_0_0_451 (.A(n_0_0_348), .B1(n_0_0_352), .B2(n_0_2), .C1(n_0_10), 
      .C2(n_0_0_353), .ZN(n_0_0_347));
   NOR2_X1 i_0_0_452 (.A1(n_0_0_368), .A2(n_0_59), .ZN(n_0_0_348));
   OAI22_X1 i_0_0_453 (.A1(n_0_106), .A2(n_0_17), .B1(n_0_18), .B2(n_0_0_403), 
      .ZN(n_0_0_349));
   AOI221_X1 i_0_0_454 (.A(n_0_0_354), .B1(n_0_0_350), .B2(n_0_0_363), .C1(
      n_0_0_355), .C2(n_0_0_364), .ZN(Sum[18]));
   MUX2_X1 i_0_0_455 (.A(n_0_0_360), .B(n_0_0_351), .S(n_0_58), .Z(n_0_0_350));
   AOI222_X1 i_0_0_456 (.A1(n_0_0_457), .A2(n_0_0_381), .B1(n_0_0_353), .B2(
      n_0_11), .C1(n_0_0_352), .C2(n_0_3), .ZN(n_0_0_351));
   NOR2_X1 i_0_0_457 (.A1(n_0_0_457), .A2(n_0_0_396), .ZN(n_0_0_352));
   NOR2_X1 i_0_0_458 (.A1(n_0_0_457), .A2(n_0_0_398), .ZN(n_0_0_353));
   OAI22_X1 i_0_0_459 (.A1(n_0_106), .A2(n_0_18), .B1(n_0_19), .B2(n_0_0_403), 
      .ZN(n_0_0_354));
   AOI221_X1 i_0_0_460 (.A(n_0_0_358), .B1(n_0_0_359), .B2(n_0_0_364), .C1(
      n_0_0_363), .C2(n_0_0_355), .ZN(Sum[19]));
   MUX2_X1 i_0_0_461 (.A(n_0_0_367), .B(n_0_0_356), .S(n_0_58), .Z(n_0_0_355));
   MUX2_X1 i_0_0_462 (.A(n_0_0_357), .B(n_0_0_395), .S(n_0_0_457), .Z(n_0_0_356));
   AOI22_X1 i_0_0_463 (.A1(n_0_12), .A2(n_0_0_399), .B1(n_0_0_397), .B2(n_0_4), 
      .ZN(n_0_0_357));
   OAI22_X1 i_0_0_464 (.A1(n_0_106), .A2(n_0_19), .B1(n_0_20), .B2(n_0_0_403), 
      .ZN(n_0_0_358));
   AOI221_X1 i_0_0_465 (.A(n_0_0_362), .B1(n_0_0_359), .B2(n_0_0_363), .C1(
      n_0_0_364), .C2(n_0_0_365), .ZN(Sum[20]));
   MUX2_X1 i_0_0_466 (.A(n_0_0_378), .B(n_0_0_360), .S(n_0_58), .Z(n_0_0_359));
   MUX2_X1 i_0_0_467 (.A(n_0_0_361), .B(n_0_0_376), .S(n_0_0_457), .Z(n_0_0_360));
   AOI22_X1 i_0_0_468 (.A1(n_0_13), .A2(n_0_0_399), .B1(n_0_0_397), .B2(n_0_5), 
      .ZN(n_0_0_361));
   OAI22_X1 i_0_0_469 (.A1(n_0_106), .A2(n_0_20), .B1(n_0_21), .B2(n_0_0_403), 
      .ZN(n_0_0_362));
   AOI221_X1 i_0_0_470 (.A(n_0_0_369), .B1(n_0_0_365), .B2(n_0_0_363), .C1(
      n_0_0_364), .C2(n_0_0_372), .ZN(Sum[21]));
   NOR2_X1 i_0_0_471 (.A1(n_0_0_404), .A2(num_leading_zeros[0]), .ZN(n_0_0_363));
   NOR2_X1 i_0_0_472 (.A1(n_0_57), .A2(n_0_0_404), .ZN(n_0_0_364));
   OAI21_X1 i_0_0_473 (.A(n_0_0_366), .B1(n_0_0_390), .B2(n_0_58), .ZN(n_0_0_365));
   NAND2_X1 i_0_0_474 (.A1(n_0_0_367), .A2(n_0_58), .ZN(n_0_0_366));
   MUX2_X1 i_0_0_475 (.A(n_0_0_368), .B(n_0_0_388), .S(n_0_0_457), .Z(n_0_0_367));
   AOI22_X1 i_0_0_476 (.A1(n_0_14), .A2(n_0_0_399), .B1(n_0_0_397), .B2(n_0_6), 
      .ZN(n_0_0_368));
   OAI22_X1 i_0_0_477 (.A1(n_0_106), .A2(n_0_21), .B1(n_0_22), .B2(n_0_0_403), 
      .ZN(n_0_0_369));
   AOI21_X1 i_0_0_478 (.A(n_0_0_402), .B1(n_0_0_370), .B2(n_0_111), .ZN(Sum[22]));
   OAI21_X1 i_0_0_479 (.A(n_0_0_383), .B1(n_0_0_371), .B2(num_leading_zeros[0]), 
      .ZN(n_0_0_370));
   INV_X1 i_0_0_480 (.A(n_0_0_372), .ZN(n_0_0_371));
   OAI21_X1 i_0_0_481 (.A(n_0_0_373), .B1(n_0_0_374), .B2(n_0_58), .ZN(n_0_0_372));
   NAND2_X1 i_0_0_482 (.A1(n_0_0_378), .A2(n_0_58), .ZN(n_0_0_373));
   OAI21_X1 i_0_0_483 (.A(n_0_0_375), .B1(n_0_0_376), .B2(n_0_0_457), .ZN(
      n_0_0_374));
   AOI222_X1 i_0_0_484 (.A1(n_0_21), .A2(n_0_0_394), .B1(n_0_0_393), .B2(n_0_5), 
      .C1(n_0_0_392), .C2(n_0_13), .ZN(n_0_0_375));
   AOI221_X1 i_0_0_485 (.A(n_0_0_377), .B1(n_0_0_397), .B2(n_0_9), .C1(n_0_17), 
      .C2(n_0_0_399), .ZN(n_0_0_376));
   NOR3_X1 i_0_0_486 (.A1(n_0_60), .A2(n_0_0_437), .A3(n_0_0_438), .ZN(n_0_0_377));
   AOI221_X1 i_0_0_487 (.A(n_0_0_379), .B1(n_0_0_394), .B2(n_0_19), .C1(n_0_59), 
      .C2(n_0_0_381), .ZN(n_0_0_378));
   INV_X1 i_0_0_488 (.A(n_0_0_380), .ZN(n_0_0_379));
   AOI22_X1 i_0_0_489 (.A1(n_0_3), .A2(n_0_0_393), .B1(n_0_0_392), .B2(n_0_11), 
      .ZN(n_0_0_380));
   INV_X1 i_0_0_490 (.A(n_0_0_382), .ZN(n_0_0_381));
   AOI22_X1 i_0_0_491 (.A1(n_0_15), .A2(n_0_0_399), .B1(n_0_0_397), .B2(n_0_7), 
      .ZN(n_0_0_382));
   OAI211_X1 i_0_0_492 (.A(num_leading_zeros[0]), .B(n_0_0_384), .C1(n_0_0_385), 
      .C2(n_0_58), .ZN(n_0_0_383));
   NAND2_X1 i_0_0_493 (.A1(n_0_58), .A2(n_0_0_390), .ZN(n_0_0_384));
   AOI21_X1 i_0_0_494 (.A(n_0_0_386), .B1(n_0_0_394), .B2(n_0_22), .ZN(n_0_0_385));
   AOI21_X1 i_0_0_495 (.A(n_0_0_387), .B1(n_0_0_388), .B2(n_0_59), .ZN(n_0_0_386));
   AOI221_X1 i_0_0_496 (.A(n_0_59), .B1(n_0_6), .B2(n_0_0_401), .C1(n_0_0_397), 
      .C2(n_0_14), .ZN(n_0_0_387));
   AOI221_X1 i_0_0_497 (.A(n_0_0_389), .B1(n_0_0_397), .B2(n_0_10), .C1(n_0_18), 
      .C2(n_0_0_399), .ZN(n_0_0_388));
   AND2_X1 i_0_0_498 (.A1(n_0_2), .A2(n_0_0_401), .ZN(n_0_0_389));
   OAI21_X1 i_0_0_499 (.A(n_0_0_391), .B1(n_0_0_395), .B2(n_0_0_457), .ZN(
      n_0_0_390));
   AOI222_X1 i_0_0_500 (.A1(n_0_20), .A2(n_0_0_394), .B1(n_0_0_393), .B2(n_0_4), 
      .C1(n_0_0_392), .C2(n_0_12), .ZN(n_0_0_391));
   NOR2_X1 i_0_0_501 (.A1(n_0_0_396), .A2(n_0_59), .ZN(n_0_0_392));
   NOR3_X1 i_0_0_502 (.A1(n_0_60), .A2(n_0_59), .A3(n_0_0_437), .ZN(n_0_0_393));
   NOR2_X1 i_0_0_503 (.A1(n_0_0_398), .A2(n_0_59), .ZN(n_0_0_394));
   AOI221_X1 i_0_0_504 (.A(n_0_0_400), .B1(n_0_0_399), .B2(n_0_16), .C1(
      n_0_0_397), .C2(n_0_8), .ZN(n_0_0_395));
   INV_X1 i_0_0_505 (.A(n_0_0_397), .ZN(n_0_0_396));
   AND2_X1 i_0_0_506 (.A1(n_0_60), .A2(n_0_0_437), .ZN(n_0_0_397));
   INV_X1 i_0_0_507 (.A(n_0_0_399), .ZN(n_0_0_398));
   NOR2_X1 i_0_0_508 (.A1(n_0_61), .A2(n_0_60), .ZN(n_0_0_399));
   AND2_X1 i_0_0_509 (.A1(n_0_0), .A2(n_0_0_401), .ZN(n_0_0_400));
   NOR2_X1 i_0_0_510 (.A1(n_0_60), .A2(n_0_0_437), .ZN(n_0_0_401));
   OAI22_X1 i_0_0_511 (.A1(n_0_106), .A2(n_0_22), .B1(n_0_23), .B2(n_0_0_403), 
      .ZN(n_0_0_402));
   NAND2_X1 i_0_0_512 (.A1(n_0_0_404), .A2(n_0_0_403), .ZN(n_0_106));
   NAND2_X1 i_0_0_513 (.A1(n_0_24), .A2(n_0_0_408), .ZN(n_0_0_403));
   INV_X1 i_0_0_514 (.A(n_0_0_404), .ZN(n_0_111));
   NAND2_X1 i_0_0_515 (.A1(n_0_0_407), .A2(n_0_0_406), .ZN(n_0_0_404));
   INV_X1 i_0_0_516 (.A(n_0_0_406), .ZN(n_0_0_405));
   NAND2_X1 i_0_0_517 (.A1(num_leading_zeros[4]), .A2(num_leading_zeros[3]), 
      .ZN(n_0_0_406));
   XNOR2_X1 i_0_0_518 (.A(B[31]), .B(n_0_0_449), .ZN(n_0_0_407));
   XNOR2_X1 i_0_0_519 (.A(B[31]), .B(A[31]), .ZN(n_0_0_408));
   OAI21_X1 i_0_0_520 (.A(n_0_0_409), .B1(n_0_0_410), .B2(n_0_0_449), .ZN(
      Sum[31]));
   NAND2_X1 i_0_0_521 (.A1(n_0_0_410), .A2(B[31]), .ZN(n_0_0_409));
   NAND2_X1 i_0_0_522 (.A1(n_0_0_413), .A2(n_0_0_411), .ZN(n_0_0_410));
   OAI21_X1 i_0_0_523 (.A(n_0_0_412), .B1(n_0_0_414), .B2(n_0_0_415), .ZN(
      n_0_0_411));
   NAND2_X1 i_0_0_524 (.A1(n_0_0_456), .A2(A[30]), .ZN(n_0_0_412));
   NAND2_X1 i_0_0_525 (.A1(n_0_0_448), .A2(B[30]), .ZN(n_0_0_413));
   AND2_X1 i_0_0_526 (.A1(n_0_0_447), .A2(B[29]), .ZN(n_0_0_414));
   AOI21_X1 i_0_0_527 (.A(n_0_0_436), .B1(n_0_0_422), .B2(n_0_0_416), .ZN(
      n_0_0_415));
   NAND2_X1 i_0_0_528 (.A1(n_0_0_419), .A2(n_0_0_417), .ZN(n_0_0_416));
   NAND2_X1 i_0_0_529 (.A1(n_0_0_455), .A2(A[28]), .ZN(n_0_0_417));
   NOR2_X1 i_0_0_530 (.A1(n_0_0_446), .A2(B[28]), .ZN(n_0_0_418));
   OAI21_X1 i_0_0_531 (.A(n_0_0_421), .B1(n_0_0_420), .B2(n_0_0_424), .ZN(
      n_0_0_419));
   NOR2_X1 i_0_0_532 (.A1(n_0_0_445), .A2(B[27]), .ZN(n_0_0_420));
   NAND2_X1 i_0_0_533 (.A1(n_0_0_445), .A2(B[27]), .ZN(n_0_0_421));
   NAND2_X1 i_0_0_534 (.A1(n_0_0_446), .A2(B[28]), .ZN(n_0_0_422));
   NOR2_X1 i_0_0_535 (.A1(n_0_0_455), .A2(A[28]), .ZN(n_0_0_423));
   AOI21_X1 i_0_0_536 (.A(n_0_0_427), .B1(n_0_0_425), .B2(n_0_0_428), .ZN(
      n_0_0_424));
   NAND2_X1 i_0_0_537 (.A1(n_0_0_454), .A2(A[26]), .ZN(n_0_0_425));
   NAND2_X1 i_0_0_538 (.A1(n_0_0_444), .A2(B[26]), .ZN(n_0_0_426));
   NOR2_X1 i_0_0_539 (.A1(n_0_0_454), .A2(A[26]), .ZN(n_0_0_427));
   OAI21_X1 i_0_0_540 (.A(n_0_0_429), .B1(n_0_0_430), .B2(n_0_0_435), .ZN(
      n_0_0_428));
   NAND2_X1 i_0_0_541 (.A1(n_0_0_443), .A2(B[25]), .ZN(n_0_0_429));
   OAI21_X1 i_0_0_542 (.A(n_0_0_431), .B1(n_0_0_432), .B2(n_0_0_433), .ZN(
      n_0_0_430));
   NAND2_X1 i_0_0_543 (.A1(n_0_0_453), .A2(A[24]), .ZN(n_0_0_431));
   NOR2_X1 i_0_0_544 (.A1(n_0_0_453), .A2(A[24]), .ZN(n_0_0_432));
   NAND2_X1 i_0_0_545 (.A1(n_0_0_452), .A2(A[23]), .ZN(n_0_0_433));
   NOR2_X1 i_0_0_546 (.A1(n_0_0_442), .A2(B[23]), .ZN(n_0_0_434));
   NOR2_X1 i_0_0_547 (.A1(n_0_0_443), .A2(B[25]), .ZN(n_0_0_435));
   NOR2_X1 i_0_0_548 (.A1(n_0_0_447), .A2(B[29]), .ZN(n_0_0_436));
   INV_X1 i_0_0_549 (.A(n_0_0_437), .ZN(n_0_61));
   XNOR2_X1 i_0_0_550 (.A(num_leading_zeros[4]), .B(n_0_0_2), .ZN(n_0_0_437));
   INV_X1 i_0_0_551 (.A(n_0_1), .ZN(n_0_0_438));
   INV_X1 i_0_0_552 (.A(num_leading_zeros[0]), .ZN(n_0_57));
   INV_X1 i_0_0_553 (.A(A[7]), .ZN(n_0_0_439));
   INV_X1 i_0_0_554 (.A(A[20]), .ZN(n_0_0_440));
   INV_X1 i_0_0_555 (.A(A[21]), .ZN(n_0_0_441));
   INV_X1 i_0_0_556 (.A(A[23]), .ZN(n_0_0_442));
   INV_X1 i_0_0_557 (.A(A[25]), .ZN(n_0_0_443));
   INV_X1 i_0_0_558 (.A(A[26]), .ZN(n_0_0_444));
   INV_X1 i_0_0_559 (.A(A[27]), .ZN(n_0_0_445));
   INV_X1 i_0_0_560 (.A(A[28]), .ZN(n_0_0_446));
   INV_X1 i_0_0_561 (.A(A[29]), .ZN(n_0_0_447));
   INV_X1 i_0_0_562 (.A(A[30]), .ZN(n_0_0_448));
   INV_X1 i_0_0_563 (.A(A[31]), .ZN(n_0_0_449));
   INV_X1 i_0_0_564 (.A(B[7]), .ZN(n_0_0_450));
   INV_X1 i_0_0_565 (.A(B[20]), .ZN(n_0_0_451));
   INV_X1 i_0_0_566 (.A(B[23]), .ZN(n_0_0_452));
   INV_X1 i_0_0_567 (.A(B[24]), .ZN(n_0_0_453));
   INV_X1 i_0_0_568 (.A(B[26]), .ZN(n_0_0_454));
   INV_X1 i_0_0_569 (.A(B[28]), .ZN(n_0_0_455));
   INV_X1 i_0_0_570 (.A(B[30]), .ZN(n_0_0_456));
   INV_X1 i_0_0_571 (.A(n_0_59), .ZN(n_0_0_457));
   INV_X1 i_0_0_572 (.A(n_0_0_410), .ZN(n_0_0_458));
   INV_X1 i_0_0_573 (.A(n_0_0_253), .ZN(n_0_0_459));
   INV_X1 i_0_0_574 (.A(n_0_0_249), .ZN(n_0_0_460));
   INV_X1 i_0_0_575 (.A(n_0_0_275), .ZN(n_0_0_461));
   INV_X1 i_0_0_576 (.A(n_0_0_124), .ZN(n_0_0_462));
endmodule
