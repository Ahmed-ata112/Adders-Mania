/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Thu Oct 27 18:49:59 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 453883483 */

module datapath(b, a, sum);
   input [31:0]b;
   input [31:0]a;
   output [32:0]sum;

   HA_X1 i_0 (.A(b[0]), .B(a[0]), .CO(n_0), .S(sum[0]));
   FA_X1 i_1 (.A(b[1]), .B(a[1]), .CI(n_0), .CO(n_1), .S(sum[1]));
   FA_X1 i_2 (.A(b[2]), .B(a[2]), .CI(n_1), .CO(n_2), .S(sum[2]));
   FA_X1 i_3 (.A(b[3]), .B(a[3]), .CI(n_2), .CO(n_3), .S(sum[3]));
   FA_X1 i_4 (.A(b[4]), .B(a[4]), .CI(n_3), .CO(n_4), .S(sum[4]));
   FA_X1 i_5 (.A(b[5]), .B(a[5]), .CI(n_4), .CO(n_5), .S(sum[5]));
   FA_X1 i_6 (.A(b[6]), .B(a[6]), .CI(n_5), .CO(n_6), .S(sum[6]));
   FA_X1 i_7 (.A(b[7]), .B(a[7]), .CI(n_6), .CO(n_7), .S(sum[7]));
   FA_X1 i_8 (.A(b[8]), .B(a[8]), .CI(n_7), .CO(n_8), .S(sum[8]));
   FA_X1 i_9 (.A(b[9]), .B(a[9]), .CI(n_8), .CO(n_9), .S(sum[9]));
   FA_X1 i_10 (.A(b[10]), .B(a[10]), .CI(n_9), .CO(n_10), .S(sum[10]));
   FA_X1 i_11 (.A(b[11]), .B(a[11]), .CI(n_10), .CO(n_11), .S(sum[11]));
   FA_X1 i_12 (.A(b[12]), .B(a[12]), .CI(n_11), .CO(n_12), .S(sum[12]));
   FA_X1 i_13 (.A(b[13]), .B(a[13]), .CI(n_12), .CO(n_13), .S(sum[13]));
   FA_X1 i_14 (.A(b[14]), .B(a[14]), .CI(n_13), .CO(n_14), .S(sum[14]));
   FA_X1 i_15 (.A(b[15]), .B(a[15]), .CI(n_14), .CO(n_15), .S(sum[15]));
   FA_X1 i_16 (.A(b[16]), .B(a[16]), .CI(n_15), .CO(n_16), .S(sum[16]));
   FA_X1 i_17 (.A(b[17]), .B(a[17]), .CI(n_16), .CO(n_17), .S(sum[17]));
   FA_X1 i_18 (.A(b[18]), .B(a[18]), .CI(n_17), .CO(n_18), .S(sum[18]));
   FA_X1 i_19 (.A(b[19]), .B(a[19]), .CI(n_18), .CO(n_19), .S(sum[19]));
   FA_X1 i_20 (.A(b[20]), .B(a[20]), .CI(n_19), .CO(n_20), .S(sum[20]));
   FA_X1 i_21 (.A(b[21]), .B(a[21]), .CI(n_20), .CO(n_21), .S(sum[21]));
   FA_X1 i_22 (.A(b[22]), .B(a[22]), .CI(n_21), .CO(n_22), .S(sum[22]));
   FA_X1 i_23 (.A(b[23]), .B(a[23]), .CI(n_22), .CO(n_23), .S(sum[23]));
   FA_X1 i_24 (.A(1'b0), .B(a[24]), .CI(n_23), .CO(n_24), .S(sum[24]));
endmodule

module simpleAdder(a, b, S, carry);
   input [31:0]a;
   input [31:0]b;
   output [31:0]S;
   output carry;

   datapath i_0 (.b({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, uc_0, b[23], 
      b[22], b[21], b[20], b[19], b[18], b[17], b[16], b[15], b[14], b[13], 
      b[12], b[11], b[10], b[9], b[8], b[7], b[6], b[5], b[4], b[3], b[2], b[1], 
      b[0]}), .a({uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, a[31], a[23], a[22], 
      a[21], a[20], a[19], a[18], a[17], a[16], a[15], a[14], a[13], a[12], 
      a[11], a[10], a[9], a[8], a[7], a[6], a[5], a[4], a[3], a[2], a[1], a[0]}), 
      .sum({uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, S[24], S[23], 
      S[22], S[21], S[20], S[19], S[18], S[17], S[16], S[15], S[14], S[13], 
      S[12], S[11], S[10], S[9], S[8], S[7], S[6], S[5], S[4], S[3], S[2], S[1], 
      S[0]}));
endmodule

module count_leading_zeros(valueIn, result);
   input [23:0]valueIn;
   output [4:0]result;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;

   AOI21_X1 i_0_0 (.A(valueIn[23]), .B1(n_0_0), .B2(n_0_9), .ZN(result[0]));
   OAI21_X1 i_0_1 (.A(n_0_1), .B1(n_0_2), .B2(valueIn[16]), .ZN(n_0_0));
   NOR3_X1 i_0_2 (.A1(valueIn[21]), .A2(valueIn[19]), .A3(valueIn[17]), .ZN(
      n_0_1));
   AOI21_X1 i_0_3 (.A(valueIn[15]), .B1(n_0_40), .B2(n_0_3), .ZN(n_0_2));
   OAI21_X1 i_0_4 (.A(n_0_39), .B1(valueIn[12]), .B2(n_0_4), .ZN(n_0_3));
   AOI21_X1 i_0_5 (.A(valueIn[11]), .B1(n_0_38), .B2(n_0_5), .ZN(n_0_4));
   OAI21_X1 i_0_6 (.A(n_0_37), .B1(valueIn[8]), .B2(n_0_6), .ZN(n_0_5));
   AOI21_X1 i_0_7 (.A(valueIn[7]), .B1(n_0_36), .B2(n_0_7), .ZN(n_0_6));
   OAI21_X1 i_0_8 (.A(n_0_35), .B1(valueIn[4]), .B2(n_0_8), .ZN(n_0_7));
   AOI21_X1 i_0_9 (.A(valueIn[3]), .B1(n_0_34), .B2(valueIn[1]), .ZN(n_0_8));
   NOR2_X1 i_0_10 (.A1(valueIn[22]), .A2(n_0_10), .ZN(n_0_9));
   NOR2_X1 i_0_11 (.A1(valueIn[21]), .A2(n_0_11), .ZN(n_0_10));
   AOI21_X1 i_0_12 (.A(valueIn[20]), .B1(n_0_41), .B2(valueIn[18]), .ZN(n_0_11));
   NOR3_X1 i_0_13 (.A1(valueIn[23]), .A2(valueIn[22]), .A3(n_0_12), .ZN(
      result[1]));
   NOR3_X1 i_0_14 (.A1(valueIn[21]), .A2(valueIn[20]), .A3(n_0_13), .ZN(n_0_12));
   NOR3_X1 i_0_15 (.A1(valueIn[19]), .A2(valueIn[18]), .A3(n_0_14), .ZN(n_0_13));
   NOR3_X1 i_0_16 (.A1(valueIn[17]), .A2(valueIn[16]), .A3(n_0_15), .ZN(n_0_14));
   NOR3_X1 i_0_17 (.A1(valueIn[15]), .A2(valueIn[14]), .A3(n_0_16), .ZN(n_0_15));
   AOI211_X1 i_0_18 (.A(valueIn[13]), .B(valueIn[12]), .C1(n_0_17), .C2(n_0_29), 
      .ZN(n_0_16));
   OAI21_X1 i_0_19 (.A(n_0_28), .B1(n_0_18), .B2(n_0_25), .ZN(n_0_17));
   NOR3_X1 i_0_20 (.A1(valueIn[5]), .A2(valueIn[4]), .A3(n_0_23), .ZN(n_0_18));
   AND2_X1 i_0_21 (.A1(n_0_19), .A2(n_0_33), .ZN(result[2]));
   NAND2_X1 i_0_22 (.A1(n_0_20), .A2(n_0_32), .ZN(n_0_19));
   OAI21_X1 i_0_23 (.A(n_0_30), .B1(n_0_24), .B2(n_0_27), .ZN(n_0_20));
   NOR2_X1 i_0_24 (.A1(n_0_21), .A2(n_0_31), .ZN(result[3]));
   AOI21_X1 i_0_25 (.A(n_0_26), .B1(n_0_24), .B2(n_0_22), .ZN(n_0_21));
   NOR4_X1 i_0_26 (.A1(valueIn[3]), .A2(valueIn[2]), .A3(valueIn[1]), .A4(
      valueIn[0]), .ZN(n_0_22));
   NOR2_X1 i_0_27 (.A1(valueIn[3]), .A2(valueIn[2]), .ZN(n_0_23));
   NOR3_X1 i_0_28 (.A1(n_0_25), .A2(valueIn[4]), .A3(valueIn[5]), .ZN(n_0_24));
   OR2_X1 i_0_29 (.A1(valueIn[7]), .A2(valueIn[6]), .ZN(n_0_25));
   NOR2_X1 i_0_30 (.A1(n_0_31), .A2(n_0_26), .ZN(result[4]));
   NAND3_X1 i_0_31 (.A1(n_0_30), .A2(n_0_29), .A3(n_0_28), .ZN(n_0_26));
   NAND2_X1 i_0_32 (.A1(n_0_29), .A2(n_0_28), .ZN(n_0_27));
   NOR2_X1 i_0_33 (.A1(valueIn[9]), .A2(valueIn[8]), .ZN(n_0_28));
   NOR2_X1 i_0_34 (.A1(valueIn[11]), .A2(valueIn[10]), .ZN(n_0_29));
   NOR4_X1 i_0_35 (.A1(valueIn[15]), .A2(valueIn[14]), .A3(valueIn[13]), 
      .A4(valueIn[12]), .ZN(n_0_30));
   NAND2_X1 i_0_36 (.A1(n_0_33), .A2(n_0_32), .ZN(n_0_31));
   NOR4_X1 i_0_37 (.A1(valueIn[19]), .A2(valueIn[18]), .A3(valueIn[17]), 
      .A4(valueIn[16]), .ZN(n_0_32));
   NOR4_X1 i_0_38 (.A1(valueIn[23]), .A2(valueIn[22]), .A3(valueIn[21]), 
      .A4(valueIn[20]), .ZN(n_0_33));
   INV_X1 i_0_39 (.A(valueIn[2]), .ZN(n_0_34));
   INV_X1 i_0_40 (.A(valueIn[5]), .ZN(n_0_35));
   INV_X1 i_0_41 (.A(valueIn[6]), .ZN(n_0_36));
   INV_X1 i_0_42 (.A(valueIn[9]), .ZN(n_0_37));
   INV_X1 i_0_43 (.A(valueIn[10]), .ZN(n_0_38));
   INV_X1 i_0_44 (.A(valueIn[13]), .ZN(n_0_39));
   INV_X1 i_0_45 (.A(valueIn[14]), .ZN(n_0_40));
   INV_X1 i_0_46 (.A(valueIn[19]), .ZN(n_0_41));
endmodule

module datapath__0_22(p_0, p_1);
   input [31:0]p_0;
   output [31:0]p_1;

   XOR2_X1 i_0 (.A(p_0[1]), .B(p_0[0]), .Z(p_1[1]));
   AND2_X1 i_1 (.A1(n_21), .A2(n_0), .ZN(p_1[2]));
   OAI21_X1 i_2 (.A(p_0[2]), .B1(p_0[1]), .B2(p_0[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(p_0[3]), .B(n_21), .Z(p_1[3]));
   XOR2_X1 i_4 (.A(p_0[4]), .B(n_20), .Z(p_1[4]));
   XOR2_X1 i_5 (.A(p_0[5]), .B(n_19), .Z(p_1[5]));
   AND2_X1 i_6 (.A1(n_18), .A2(n_1), .ZN(p_1[6]));
   OAI21_X1 i_7 (.A(p_0[6]), .B1(n_19), .B2(p_0[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(p_0[7]), .B(n_18), .Z(p_1[7]));
   XOR2_X1 i_9 (.A(p_0[8]), .B(n_17), .Z(p_1[8]));
   AND2_X1 i_10 (.A1(n_16), .A2(n_2), .ZN(p_1[9]));
   OAI21_X1 i_11 (.A(p_0[9]), .B1(n_17), .B2(p_0[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(p_0[10]), .B(n_16), .Z(p_1[10]));
   XNOR2_X1 i_13 (.A(p_0[11]), .B(n_15), .ZN(p_1[11]));
   XOR2_X1 i_14 (.A(p_0[12]), .B(n_14), .Z(p_1[12]));
   XOR2_X1 i_15 (.A(p_0[13]), .B(n_13), .Z(p_1[13]));
   XNOR2_X1 i_16 (.A(p_0[14]), .B(n_12), .ZN(p_1[14]));
   XNOR2_X1 i_17 (.A(p_0[15]), .B(n_11), .ZN(p_1[15]));
   XOR2_X1 i_18 (.A(p_0[16]), .B(n_10), .Z(p_1[16]));
   XOR2_X1 i_19 (.A(p_0[17]), .B(n_9), .Z(p_1[17]));
   XOR2_X1 i_20 (.A(p_0[18]), .B(n_8), .Z(p_1[18]));
   AND2_X1 i_21 (.A1(n_7), .A2(n_3), .ZN(p_1[19]));
   OAI21_X1 i_22 (.A(p_0[19]), .B1(n_8), .B2(p_0[18]), .ZN(n_3));
   XOR2_X1 i_23 (.A(p_0[20]), .B(n_7), .Z(p_1[20]));
   AND2_X1 i_24 (.A1(n_6), .A2(n_4), .ZN(p_1[21]));
   OAI21_X1 i_25 (.A(p_0[21]), .B1(n_7), .B2(p_0[20]), .ZN(n_4));
   XOR2_X1 i_26 (.A(p_0[22]), .B(n_6), .Z(p_1[22]));
   AND2_X1 i_27 (.A1(p_1[31]), .A2(n_5), .ZN(p_1[23]));
   OAI21_X1 i_28 (.A(p_0[23]), .B1(n_6), .B2(p_0[22]), .ZN(n_5));
   OR3_X1 i_29 (.A1(n_6), .A2(p_0[22]), .A3(p_0[23]), .ZN(p_1[31]));
   OR3_X1 i_30 (.A1(n_7), .A2(p_0[20]), .A3(p_0[21]), .ZN(n_6));
   OR3_X1 i_31 (.A1(n_8), .A2(p_0[18]), .A3(p_0[19]), .ZN(n_7));
   OR2_X1 i_32 (.A1(n_9), .A2(p_0[17]), .ZN(n_8));
   OR2_X1 i_33 (.A1(n_10), .A2(p_0[16]), .ZN(n_9));
   NAND2_X1 i_34 (.A1(n_11), .A2(n_23), .ZN(n_10));
   NOR3_X1 i_35 (.A1(n_13), .A2(p_0[13]), .A3(p_0[14]), .ZN(n_11));
   NOR2_X1 i_36 (.A1(n_13), .A2(p_0[13]), .ZN(n_12));
   OR2_X1 i_37 (.A1(n_14), .A2(p_0[12]), .ZN(n_13));
   NAND2_X1 i_38 (.A1(n_15), .A2(n_22), .ZN(n_14));
   NOR2_X1 i_39 (.A1(n_16), .A2(p_0[10]), .ZN(n_15));
   OR3_X1 i_40 (.A1(n_17), .A2(p_0[8]), .A3(p_0[9]), .ZN(n_16));
   OR2_X1 i_41 (.A1(n_18), .A2(p_0[7]), .ZN(n_17));
   OR3_X1 i_42 (.A1(n_19), .A2(p_0[5]), .A3(p_0[6]), .ZN(n_18));
   OR2_X1 i_43 (.A1(n_20), .A2(p_0[4]), .ZN(n_19));
   OR2_X1 i_44 (.A1(n_21), .A2(p_0[3]), .ZN(n_20));
   OR3_X1 i_45 (.A1(p_0[2]), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_21));
   INV_X1 i_46 (.A(p_0[11]), .ZN(n_22));
   INV_X1 i_47 (.A(p_0[15]), .ZN(n_23));
endmodule

module fp_adder(A, B, Sum);
   input [31:0]A;
   input [31:0]B;
   output [31:0]Sum;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire [4:0]num_leading_zeros;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire [7:0]exp_Sum;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire [31:0]mant_A_reg;
   wire n_0_49;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_50;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_51;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_52;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_53;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_54;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_55;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_56;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_57;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_58;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_59;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_60;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_61;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_62;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_63;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_64;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_65;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_66;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_67;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_68;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_69;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_70;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_71;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_72;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_73;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_74;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_75;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_76;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_77;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_78;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_79;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_80;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_81;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_82;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_83;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_84;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_85;
   wire n_0_0_231;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_86;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_87;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_88;
   wire n_0_0_246;
   wire n_0_0_247;
   wire n_0_0_248;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_89;
   wire n_0_0_253;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_90;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_91;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_0_266;
   wire n_0_92;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_93;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_94;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_95;
   wire n_0_0_288;
   wire n_0_0_289;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_0_304;
   wire n_0_0_305;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_0_311;
   wire n_0_0_312;
   wire n_0_0_313;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_0_321;
   wire n_0_0_322;
   wire n_0_0_323;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_328;
   wire n_0_0_329;
   wire n_0_0_330;
   wire n_0_0_331;
   wire n_0_0_332;
   wire n_0_0_333;
   wire n_0_0_334;
   wire n_0_0_335;
   wire n_0_0_336;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_341;
   wire n_0_0_342;
   wire n_0_0_343;
   wire n_0_0_344;
   wire n_0_0_345;
   wire n_0_0_346;
   wire n_0_0_347;
   wire n_0_0_348;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_351;
   wire n_0_0_352;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_0_355;
   wire n_0_0_356;
   wire n_0_0_357;
   wire n_0_0_358;
   wire n_0_0_359;
   wire n_0_0_360;
   wire n_0_0_361;
   wire n_0_0_362;
   wire n_0_0_363;
   wire n_0_0_364;
   wire n_0_0_365;
   wire n_0_0_366;
   wire n_0_0_367;
   wire n_0_0_368;
   wire n_0_0_369;
   wire n_0_0_370;
   wire n_0_0_371;
   wire n_0_0_372;
   wire n_0_0_373;
   wire n_0_0_374;
   wire n_0_0_375;
   wire n_0_0_376;
   wire n_0_0_377;
   wire n_0_0_378;
   wire n_0_0_379;
   wire n_0_0_380;
   wire n_0_0_381;
   wire n_0_0_382;
   wire n_0_0_383;
   wire n_0_0_384;
   wire n_0_0_385;
   wire n_0_0_386;
   wire n_0_0_387;
   wire n_0_0_388;
   wire n_0_0_389;
   wire n_0_0_390;
   wire n_0_0_391;
   wire n_0_0_392;
   wire n_0_0_393;
   wire n_0_0_394;
   wire n_0_0_395;
   wire n_0_0_396;
   wire n_0_0_397;
   wire n_0_0_398;
   wire n_0_0_399;
   wire n_0_0_400;
   wire n_0_0_401;
   wire n_0_0_402;
   wire n_0_0_403;
   wire n_0_0_404;
   wire n_0_0_405;
   wire n_0_0_406;
   wire n_0_0_407;
   wire n_0_0_408;
   wire n_0_0_409;
   wire n_0_0_410;
   wire n_0_0_411;
   wire n_0_0_412;
   wire n_0_0_413;
   wire n_0_0_414;
   wire n_0_0_415;
   wire n_0_0_416;
   wire n_0_0_417;
   wire n_0_0_418;
   wire n_0_0_419;
   wire n_0_0_420;
   wire n_0_0_421;
   wire n_0_0_422;
   wire n_0_0_423;
   wire n_0_0_424;
   wire n_0_0_425;
   wire n_0_0_426;
   wire n_0_0_427;
   wire n_0_0_428;
   wire n_0_0_429;
   wire n_0_0_430;
   wire n_0_0_431;
   wire n_0_0_432;
   wire n_0_0_433;
   wire n_0_0_434;
   wire n_0_0_435;
   wire n_0_0_436;
   wire n_0_0_437;
   wire n_0_0_438;
   wire n_0_0_439;
   wire n_0_0_440;
   wire n_0_0_441;
   wire n_0_0_442;
   wire n_0_0_443;
   wire n_0_0_444;
   wire n_0_0_445;
   wire n_0_0_446;
   wire n_0_0_447;
   wire n_0_0_448;
   wire n_0_0_449;
   wire n_0_0_450;
   wire n_0_0_451;
   wire n_0_0_452;
   wire n_0_0_453;
   wire n_0_0_454;
   wire n_0_0_455;
   wire n_0_0_456;
   wire n_0_0_457;
   wire n_0_0_458;
   wire n_0_0_459;
   wire n_0_0_460;
   wire n_0_0_461;
   wire n_0_0_462;
   wire n_0_0_463;
   wire n_0_0_464;
   wire n_0_0_465;
   wire n_0_0_466;
   wire n_0_0_467;
   wire n_0_0_468;
   wire n_0_0_469;
   wire n_0_0_470;
   wire n_0_0_471;
   wire n_0_0_472;
   wire n_0_0_473;
   wire n_0_96;
   wire n_0_0_474;
   wire n_0_0_475;
   wire n_0_0_476;
   wire n_0_0_477;
   wire n_0_0_478;
   wire n_0_0_479;
   wire n_0_0_480;
   wire n_0_0_481;
   wire n_0_0_482;
   wire n_0_0_483;
   wire n_0_0_484;
   wire n_0_0_485;
   wire n_0_0_486;
   wire n_0_0_487;
   wire n_0_0_488;
   wire n_0_0_489;
   wire n_0_0_490;
   wire n_0_0_491;
   wire n_0_0_492;
   wire n_0_0_493;
   wire n_0_0_494;
   wire n_0_0_495;
   wire n_0_0_496;
   wire n_0_0_497;
   wire n_0_0_498;
   wire n_0_0_499;
   wire n_0_0_500;
   wire n_0_0_501;
   wire n_0_0_502;
   wire n_0_0_503;
   wire n_0_0_504;
   wire n_0_0_505;
   wire n_0_0_506;
   wire n_0_0_507;
   wire n_0_0_508;
   wire n_0_0_509;
   wire n_0_0_510;
   wire n_0_0_511;
   wire n_0_0_512;
   wire n_0_0_513;
   wire n_0_0_514;
   wire n_0_0_515;
   wire n_0_0_516;
   wire n_0_0_517;
   wire n_0_0_518;
   wire n_0_0_519;
   wire n_0_0_520;
   wire n_0_0_521;
   wire n_0_0_522;
   wire n_0_0_523;
   wire n_0_0_524;
   wire n_0_0_525;
   wire n_0_0_526;
   wire n_0_0_527;

   simpleAdder simpleAdder_dut (.a({mant_A_reg[31], uc_0, uc_1, uc_2, uc_3, uc_4, 
      uc_5, uc_6, mant_A_reg[23], mant_A_reg[22], mant_A_reg[21], mant_A_reg[20], 
      mant_A_reg[19], mant_A_reg[18], mant_A_reg[17], mant_A_reg[16], 
      mant_A_reg[15], mant_A_reg[14], mant_A_reg[13], mant_A_reg[12], 
      mant_A_reg[11], mant_A_reg[10], mant_A_reg[9], mant_A_reg[8], 
      mant_A_reg[7], mant_A_reg[6], mant_A_reg[5], mant_A_reg[4], mant_A_reg[3], 
      mant_A_reg[2], mant_A_reg[1], n_0_49}), .b({uc_7, uc_8, uc_9, uc_10, uc_11, 
      uc_12, uc_13, uc_14, n_0_96, n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, 
      n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, 
      n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73}), 
      .S({uc_15, uc_16, uc_17, uc_18, uc_19, uc_20, uc_21, n_0_24, n_0_23, 
      n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, 
      n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, 
      n_0_3, n_0_2, n_0_1, n_0_0}), .carry());
   count_leading_zeros count_leading_zeros_instance (.valueIn({n_0_23, n_0_22, 
      n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, 
      n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, 
      n_0_2, n_0_1, n_0_0}), .result(num_leading_zeros));
   datapath__0_22 i_0_14 (.p_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, 
      n_0_63, n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, 
      n_0_54, n_0_53, n_0_52, n_0_51, n_0_50, n_0_49}), .p_1({n_0_48, uc_22, 
      uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, n_0_47, n_0_46, n_0_45, n_0_44, 
      n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, 
      n_0_34, n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, 
      n_0_25, uc_29}));
   HA_X1 i_0_0_0 (.A(n_0_24), .B(n_0_0_462), .CO(n_0_0_0), .S(exp_Sum[0]));
   HA_X1 i_0_0_1 (.A(n_0_0_464), .B(n_0_0_0), .CO(n_0_0_1), .S(exp_Sum[1]));
   HA_X1 i_0_0_2 (.A(n_0_0_455), .B(n_0_0_1), .CO(n_0_0_2), .S(exp_Sum[2]));
   HA_X1 i_0_0_3 (.A(n_0_0_466), .B(n_0_0_2), .CO(n_0_0_3), .S(exp_Sum[3]));
   HA_X1 i_0_0_4 (.A(n_0_0_471), .B(n_0_0_3), .CO(n_0_0_4), .S(exp_Sum[4]));
   HA_X1 i_0_0_5 (.A(n_0_0_445), .B(n_0_0_4), .CO(n_0_0_5), .S(exp_Sum[5]));
   HA_X1 i_0_0_6 (.A(n_0_0_440), .B(n_0_0_5), .CO(n_0_0_6), .S(exp_Sum[6]));
   MUX2_X1 i_0_0_7 (.A(n_0_25), .B(n_0_50), .S(n_0_0_442), .Z(mant_A_reg[1]));
   MUX2_X1 i_0_0_8 (.A(n_0_26), .B(n_0_51), .S(n_0_0_442), .Z(mant_A_reg[2]));
   MUX2_X1 i_0_0_9 (.A(n_0_27), .B(n_0_52), .S(n_0_0_442), .Z(mant_A_reg[3]));
   MUX2_X1 i_0_0_10 (.A(n_0_28), .B(n_0_53), .S(n_0_0_442), .Z(mant_A_reg[4]));
   MUX2_X1 i_0_0_11 (.A(n_0_29), .B(n_0_54), .S(n_0_0_442), .Z(mant_A_reg[5]));
   MUX2_X1 i_0_0_12 (.A(n_0_30), .B(n_0_55), .S(n_0_0_442), .Z(mant_A_reg[6]));
   MUX2_X1 i_0_0_13 (.A(n_0_31), .B(n_0_56), .S(n_0_0_442), .Z(mant_A_reg[7]));
   MUX2_X1 i_0_0_14 (.A(n_0_32), .B(n_0_57), .S(n_0_0_442), .Z(mant_A_reg[8]));
   MUX2_X1 i_0_0_15 (.A(n_0_33), .B(n_0_58), .S(n_0_0_442), .Z(mant_A_reg[9]));
   MUX2_X1 i_0_0_16 (.A(n_0_34), .B(n_0_59), .S(n_0_0_442), .Z(mant_A_reg[10]));
   MUX2_X1 i_0_0_17 (.A(n_0_35), .B(n_0_60), .S(n_0_0_442), .Z(mant_A_reg[11]));
   MUX2_X1 i_0_0_18 (.A(n_0_36), .B(n_0_61), .S(n_0_0_442), .Z(mant_A_reg[12]));
   MUX2_X1 i_0_0_19 (.A(n_0_37), .B(n_0_62), .S(n_0_0_442), .Z(mant_A_reg[13]));
   MUX2_X1 i_0_0_20 (.A(n_0_38), .B(n_0_63), .S(n_0_0_442), .Z(mant_A_reg[14]));
   MUX2_X1 i_0_0_21 (.A(n_0_39), .B(n_0_64), .S(n_0_0_442), .Z(mant_A_reg[15]));
   MUX2_X1 i_0_0_22 (.A(n_0_40), .B(n_0_65), .S(n_0_0_442), .Z(mant_A_reg[16]));
   MUX2_X1 i_0_0_23 (.A(n_0_41), .B(n_0_66), .S(n_0_0_442), .Z(mant_A_reg[17]));
   MUX2_X1 i_0_0_24 (.A(n_0_42), .B(n_0_67), .S(n_0_0_442), .Z(mant_A_reg[18]));
   MUX2_X1 i_0_0_25 (.A(n_0_43), .B(n_0_68), .S(n_0_0_442), .Z(mant_A_reg[19]));
   MUX2_X1 i_0_0_26 (.A(n_0_44), .B(n_0_69), .S(n_0_0_442), .Z(mant_A_reg[20]));
   MUX2_X1 i_0_0_27 (.A(n_0_45), .B(n_0_70), .S(n_0_0_442), .Z(mant_A_reg[21]));
   MUX2_X1 i_0_0_28 (.A(n_0_46), .B(n_0_71), .S(n_0_0_442), .Z(mant_A_reg[22]));
   MUX2_X1 i_0_0_29 (.A(n_0_47), .B(n_0_72), .S(n_0_0_442), .Z(mant_A_reg[23]));
   AND2_X1 i_0_0_30 (.A1(n_0_0_520), .A2(n_0_48), .ZN(mant_A_reg[31]));
   OAI211_X1 i_0_0_31 (.A(n_0_0_8), .B(n_0_0_7), .C1(n_0_0_101), .C2(n_0_0_27), 
      .ZN(n_0_49));
   NAND2_X1 i_0_0_32 (.A1(A[0]), .A2(n_0_0_474), .ZN(n_0_0_7));
   NAND3_X1 i_0_0_33 (.A1(n_0_0_10), .A2(n_0_0_9), .A3(n_0_0_141), .ZN(n_0_0_8));
   AOI22_X1 i_0_0_34 (.A1(n_0_0_148), .A2(n_0_0_62), .B1(n_0_0_38), .B2(n_0_0_30), 
      .ZN(n_0_0_9));
   NAND2_X1 i_0_0_35 (.A1(n_0_0_12), .A2(n_0_0_11), .ZN(n_0_0_10));
   AOI21_X1 i_0_0_36 (.A(n_0_0_143), .B1(n_0_0_121), .B2(A[3]), .ZN(n_0_0_11));
   AOI222_X1 i_0_0_37 (.A1(A[0]), .A2(n_0_0_521), .B1(n_0_0_136), .B2(A[1]), 
      .C1(A[2]), .C2(n_0_0_122), .ZN(n_0_0_12));
   OAI211_X1 i_0_0_38 (.A(n_0_0_14), .B(n_0_0_13), .C1(n_0_0_107), .C2(n_0_0_27), 
      .ZN(n_0_50));
   NAND2_X1 i_0_0_39 (.A1(A[1]), .A2(n_0_0_474), .ZN(n_0_0_13));
   NAND4_X1 i_0_0_40 (.A1(n_0_0_18), .A2(n_0_0_141), .A3(n_0_0_19), .A4(n_0_0_15), 
      .ZN(n_0_0_14));
   NAND2_X1 i_0_0_41 (.A1(n_0_0_17), .A2(n_0_0_16), .ZN(n_0_0_15));
   AOI21_X1 i_0_0_42 (.A(n_0_0_143), .B1(n_0_0_123), .B2(n_0_0_34), .ZN(n_0_0_16));
   AOI222_X1 i_0_0_43 (.A1(A[1]), .A2(n_0_0_521), .B1(n_0_0_136), .B2(A[2]), 
      .C1(A[4]), .C2(n_0_0_121), .ZN(n_0_0_17));
   NAND2_X1 i_0_0_44 (.A1(n_0_0_41), .A2(n_0_0_30), .ZN(n_0_0_18));
   NAND2_X1 i_0_0_45 (.A1(n_0_0_148), .A2(n_0_0_66), .ZN(n_0_0_19));
   AOI21_X1 i_0_0_46 (.A(n_0_0_20), .B1(n_0_0_474), .B2(n_0_0_498), .ZN(n_0_51));
   AOI211_X1 i_0_0_47 (.A(n_0_0_474), .B(n_0_0_22), .C1(n_0_0_21), .C2(n_0_0_156), 
      .ZN(n_0_0_20));
   NOR2_X1 i_0_0_48 (.A1(n_0_0_148), .A2(n_0_0_113), .ZN(n_0_0_21));
   AOI211_X1 i_0_0_49 (.A(n_0_0_156), .B(n_0_0_23), .C1(n_0_0_70), .C2(n_0_0_148), 
      .ZN(n_0_0_22));
   AOI21_X1 i_0_0_50 (.A(n_0_0_148), .B1(n_0_0_25), .B2(n_0_0_24), .ZN(n_0_0_23));
   OAI211_X1 i_0_0_51 (.A(n_0_0_26), .B(n_0_0_146), .C1(n_0_0_149), .C2(
      n_0_0_498), .ZN(n_0_0_24));
   NAND2_X1 i_0_0_52 (.A1(n_0_0_145), .A2(n_0_0_52), .ZN(n_0_0_25));
   AOI22_X1 i_0_0_53 (.A1(A[3]), .A2(n_0_0_136), .B1(n_0_0_123), .B2(n_0_0_39), 
      .ZN(n_0_0_26));
   OAI211_X1 i_0_0_54 (.A(n_0_0_35), .B(n_0_0_28), .C1(n_0_0_27), .C2(n_0_0_118), 
      .ZN(n_0_52));
   NAND3_X1 i_0_0_55 (.A1(n_0_96), .A2(n_0_0_156), .A3(n_0_0_147), .ZN(n_0_0_27));
   OAI211_X1 i_0_0_56 (.A(n_0_0_141), .B(n_0_0_29), .C1(n_0_0_74), .C2(n_0_0_147), 
      .ZN(n_0_0_28));
   OAI211_X1 i_0_0_57 (.A(n_0_0_147), .B(n_0_0_31), .C1(n_0_0_56), .C2(n_0_0_146), 
      .ZN(n_0_0_29));
   NOR2_X1 i_0_0_58 (.A1(n_0_0_148), .A2(n_0_0_146), .ZN(n_0_0_30));
   NAND3_X1 i_0_0_59 (.A1(n_0_0_152), .A2(n_0_0_146), .A3(n_0_0_32), .ZN(
      n_0_0_31));
   AOI21_X1 i_0_0_60 (.A(n_0_0_33), .B1(n_0_0_43), .B2(n_0_0_151), .ZN(n_0_0_32));
   AOI211_X1 i_0_0_61 (.A(n_0_0_151), .B(n_0_0_34), .C1(A[4]), .C2(n_0_0_315), 
      .ZN(n_0_0_33));
   AND2_X1 i_0_0_62 (.A1(A[3]), .A2(n_0_0_316), .ZN(n_0_0_34));
   NAND2_X1 i_0_0_63 (.A1(A[3]), .A2(n_0_0_474), .ZN(n_0_0_35));
   OAI221_X1 i_0_0_64 (.A(n_0_0_36), .B1(n_0_0_82), .B2(n_0_0_95), .C1(n_0_0_138), 
      .C2(n_0_0_38), .ZN(n_0_53));
   INV_X1 i_0_0_65 (.A(n_0_0_37), .ZN(n_0_0_36));
   OAI221_X1 i_0_0_66 (.A(n_0_0_40), .B1(n_0_0_47), .B2(n_0_0_127), .C1(n_0_0_55), 
      .C2(n_0_0_63), .ZN(n_0_0_37));
   AOI22_X1 i_0_0_67 (.A1(n_0_0_150), .A2(n_0_0_39), .B1(n_0_0_123), .B2(
      n_0_0_53), .ZN(n_0_0_38));
   MUX2_X1 i_0_0_68 (.A(A[5]), .B(A[4]), .S(n_0_0_316), .Z(n_0_0_39));
   NAND2_X1 i_0_0_69 (.A1(A[4]), .A2(n_0_0_474), .ZN(n_0_0_40));
   OAI221_X1 i_0_0_70 (.A(n_0_0_45), .B1(n_0_0_41), .B2(n_0_0_138), .C1(n_0_0_67), 
      .C2(n_0_0_55), .ZN(n_0_54));
   AOI221_X1 i_0_0_71 (.A(n_0_0_42), .B1(n_0_0_57), .B2(n_0_0_123), .C1(A[5]), 
      .C2(n_0_0_521), .ZN(n_0_0_41));
   AND2_X1 i_0_0_72 (.A1(A[6]), .A2(n_0_0_136), .ZN(n_0_0_42));
   AOI21_X1 i_0_0_73 (.A(n_0_0_44), .B1(n_0_0_315), .B2(A[6]), .ZN(n_0_0_43));
   AND2_X1 i_0_0_74 (.A1(A[5]), .A2(n_0_0_316), .ZN(n_0_0_44));
   AOI211_X1 i_0_0_75 (.A(n_0_0_48), .B(n_0_0_46), .C1(A[5]), .C2(n_0_0_474), 
      .ZN(n_0_0_45));
   NOR2_X1 i_0_0_76 (.A1(n_0_0_130), .A2(n_0_0_47), .ZN(n_0_0_46));
   NAND3_X1 i_0_0_77 (.A1(n_0_96), .A2(n_0_0_156), .A3(n_0_0_144), .ZN(n_0_0_47));
   NOR2_X1 i_0_0_78 (.A1(n_0_0_95), .A2(n_0_0_86), .ZN(n_0_0_48));
   AOI221_X1 i_0_0_79 (.A(n_0_0_49), .B1(n_0_0_51), .B2(n_0_0_139), .C1(n_0_0_90), 
      .C2(n_0_0_96), .ZN(n_0_55));
   OAI21_X1 i_0_0_80 (.A(n_0_0_50), .B1(n_0_96), .B2(A[6]), .ZN(n_0_0_49));
   OAI211_X1 i_0_0_81 (.A(n_0_96), .B(n_0_0_156), .C1(n_0_0_135), .C2(n_0_0_143), 
      .ZN(n_0_0_50));
   MUX2_X1 i_0_0_82 (.A(n_0_0_71), .B(n_0_0_52), .S(n_0_0_146), .Z(n_0_0_51));
   AOI22_X1 i_0_0_83 (.A1(n_0_0_150), .A2(n_0_0_53), .B1(n_0_0_123), .B2(
      n_0_0_64), .ZN(n_0_0_52));
   MUX2_X1 i_0_0_84 (.A(A[7]), .B(A[6]), .S(n_0_0_316), .Z(n_0_0_53));
   AOI221_X1 i_0_0_85 (.A(n_0_0_54), .B1(n_0_0_56), .B2(n_0_0_137), .C1(n_0_0_97), 
      .C2(n_0_0_96), .ZN(n_0_56));
   OAI22_X1 i_0_0_86 (.A1(n_0_0_76), .A2(n_0_0_55), .B1(n_0_0_60), .B2(n_0_0_61), 
      .ZN(n_0_0_54));
   NAND2_X1 i_0_0_87 (.A1(n_0_0_145), .A2(n_0_0_139), .ZN(n_0_0_55));
   AOI22_X1 i_0_0_88 (.A1(n_0_0_150), .A2(n_0_0_57), .B1(n_0_0_123), .B2(
      n_0_0_68), .ZN(n_0_0_56));
   INV_X1 i_0_0_89 (.A(n_0_0_58), .ZN(n_0_0_57));
   AOI21_X1 i_0_0_90 (.A(n_0_0_59), .B1(n_0_0_315), .B2(A[8]), .ZN(n_0_0_58));
   AND2_X1 i_0_0_91 (.A1(A[7]), .A2(n_0_0_316), .ZN(n_0_0_59));
   AOI21_X1 i_0_0_92 (.A(n_0_0_474), .B1(n_0_0_156), .B2(n_0_0_142), .ZN(
      n_0_0_60));
   AND2_X1 i_0_0_93 (.A1(A[7]), .A2(n_0_0_474), .ZN(n_0_0_61));
   OAI221_X1 i_0_0_94 (.A(n_0_0_65), .B1(n_0_0_62), .B2(n_0_0_140), .C1(
      n_0_0_101), .C2(n_0_0_95), .ZN(n_0_57));
   MUX2_X1 i_0_0_95 (.A(n_0_0_83), .B(n_0_0_63), .S(n_0_0_146), .Z(n_0_0_62));
   AOI22_X1 i_0_0_96 (.A1(n_0_0_150), .A2(n_0_0_64), .B1(n_0_0_123), .B2(
      n_0_0_72), .ZN(n_0_0_63));
   MUX2_X1 i_0_0_97 (.A(A[9]), .B(A[8]), .S(n_0_0_316), .Z(n_0_0_64));
   NAND2_X1 i_0_0_98 (.A1(A[8]), .A2(n_0_0_474), .ZN(n_0_0_65));
   OAI221_X1 i_0_0_99 (.A(n_0_0_69), .B1(n_0_0_66), .B2(n_0_0_140), .C1(
      n_0_0_107), .C2(n_0_0_95), .ZN(n_0_58));
   MUX2_X1 i_0_0_100 (.A(n_0_0_87), .B(n_0_0_67), .S(n_0_0_146), .Z(n_0_0_66));
   AOI22_X1 i_0_0_101 (.A1(n_0_0_150), .A2(n_0_0_68), .B1(n_0_0_123), .B2(
      n_0_0_78), .ZN(n_0_0_67));
   MUX2_X1 i_0_0_102 (.A(A[10]), .B(A[9]), .S(n_0_0_316), .Z(n_0_0_68));
   NAND2_X1 i_0_0_103 (.A1(A[9]), .A2(n_0_0_474), .ZN(n_0_0_69));
   OAI221_X1 i_0_0_104 (.A(n_0_0_73), .B1(n_0_0_70), .B2(n_0_0_140), .C1(
      n_0_0_113), .C2(n_0_0_95), .ZN(n_0_59));
   MUX2_X1 i_0_0_105 (.A(n_0_0_91), .B(n_0_0_71), .S(n_0_0_146), .Z(n_0_0_70));
   AOI22_X1 i_0_0_106 (.A1(n_0_0_150), .A2(n_0_0_72), .B1(n_0_0_123), .B2(
      n_0_0_84), .ZN(n_0_0_71));
   MUX2_X1 i_0_0_107 (.A(A[11]), .B(A[10]), .S(n_0_0_316), .Z(n_0_0_72));
   NAND2_X1 i_0_0_108 (.A1(A[10]), .A2(n_0_0_474), .ZN(n_0_0_73));
   OAI221_X1 i_0_0_109 (.A(n_0_0_80), .B1(n_0_0_75), .B2(n_0_0_140), .C1(
      n_0_0_118), .C2(n_0_0_95), .ZN(n_0_60));
   INV_X1 i_0_0_110 (.A(n_0_0_75), .ZN(n_0_0_74));
   OAI21_X1 i_0_0_111 (.A(n_0_0_79), .B1(n_0_0_76), .B2(n_0_0_145), .ZN(n_0_0_75));
   INV_X1 i_0_0_112 (.A(n_0_0_77), .ZN(n_0_0_76));
   AOI22_X1 i_0_0_113 (.A1(n_0_0_150), .A2(n_0_0_78), .B1(n_0_0_123), .B2(
      n_0_0_88), .ZN(n_0_0_77));
   MUX2_X1 i_0_0_114 (.A(A[12]), .B(A[11]), .S(n_0_0_316), .Z(n_0_0_78));
   NAND2_X1 i_0_0_115 (.A1(n_0_0_145), .A2(n_0_0_98), .ZN(n_0_0_79));
   NAND2_X1 i_0_0_116 (.A1(A[11]), .A2(n_0_0_474), .ZN(n_0_0_80));
   OAI221_X1 i_0_0_117 (.A(n_0_0_81), .B1(n_0_0_94), .B2(n_0_0_127), .C1(
      n_0_0_140), .C2(n_0_0_82), .ZN(n_0_61));
   NAND2_X1 i_0_0_118 (.A1(A[12]), .A2(n_0_0_474), .ZN(n_0_0_81));
   MUX2_X1 i_0_0_119 (.A(n_0_0_83), .B(n_0_0_102), .S(n_0_0_145), .Z(n_0_0_82));
   AOI22_X1 i_0_0_120 (.A1(n_0_0_150), .A2(n_0_0_84), .B1(n_0_0_123), .B2(
      n_0_0_92), .ZN(n_0_0_83));
   MUX2_X1 i_0_0_121 (.A(A[13]), .B(A[12]), .S(n_0_0_316), .Z(n_0_0_84));
   OAI221_X1 i_0_0_122 (.A(n_0_0_85), .B1(n_0_0_94), .B2(n_0_0_130), .C1(
      n_0_0_140), .C2(n_0_0_86), .ZN(n_0_62));
   NAND2_X1 i_0_0_123 (.A1(A[13]), .A2(n_0_0_474), .ZN(n_0_0_85));
   MUX2_X1 i_0_0_124 (.A(n_0_0_87), .B(n_0_0_108), .S(n_0_0_145), .Z(n_0_0_86));
   AOI22_X1 i_0_0_125 (.A1(n_0_0_150), .A2(n_0_0_88), .B1(n_0_0_123), .B2(
      n_0_0_99), .ZN(n_0_0_87));
   MUX2_X1 i_0_0_126 (.A(A[14]), .B(A[13]), .S(n_0_0_316), .Z(n_0_0_88));
   OAI221_X1 i_0_0_127 (.A(n_0_0_89), .B1(n_0_0_135), .B2(n_0_0_94), .C1(
      n_0_0_90), .C2(n_0_0_140), .ZN(n_0_63));
   NAND2_X1 i_0_0_128 (.A1(A[14]), .A2(n_0_0_474), .ZN(n_0_0_89));
   MUX2_X1 i_0_0_129 (.A(n_0_0_91), .B(n_0_0_114), .S(n_0_0_145), .Z(n_0_0_90));
   AOI22_X1 i_0_0_130 (.A1(n_0_0_150), .A2(n_0_0_92), .B1(n_0_0_123), .B2(
      n_0_0_105), .ZN(n_0_0_91));
   MUX2_X1 i_0_0_131 (.A(A[15]), .B(A[14]), .S(n_0_0_316), .Z(n_0_0_92));
   OAI221_X1 i_0_0_132 (.A(n_0_0_93), .B1(n_0_0_97), .B2(n_0_0_140), .C1(
      n_0_0_149), .C2(n_0_0_94), .ZN(n_0_64));
   NAND2_X1 i_0_0_133 (.A1(A[15]), .A2(n_0_0_474), .ZN(n_0_0_93));
   NAND2_X1 i_0_0_134 (.A1(n_0_0_96), .A2(n_0_0_146), .ZN(n_0_0_94));
   NAND2_X1 i_0_0_135 (.A1(n_0_0_141), .A2(n_0_0_148), .ZN(n_0_0_95));
   NOR3_X1 i_0_0_136 (.A1(n_0_0_474), .A2(n_0_0_156), .A3(n_0_0_147), .ZN(
      n_0_0_96));
   MUX2_X1 i_0_0_137 (.A(n_0_0_98), .B(n_0_0_120), .S(n_0_0_145), .Z(n_0_0_97));
   AOI22_X1 i_0_0_138 (.A1(n_0_0_150), .A2(n_0_0_99), .B1(n_0_0_123), .B2(
      n_0_0_111), .ZN(n_0_0_98));
   MUX2_X1 i_0_0_139 (.A(A[16]), .B(A[15]), .S(n_0_0_316), .Z(n_0_0_99));
   OAI21_X1 i_0_0_140 (.A(n_0_0_100), .B1(n_0_0_101), .B2(n_0_0_140), .ZN(n_0_65));
   NAND2_X1 i_0_0_141 (.A1(A[16]), .A2(n_0_0_474), .ZN(n_0_0_100));
   MUX2_X1 i_0_0_142 (.A(n_0_0_127), .B(n_0_0_102), .S(n_0_0_146), .Z(n_0_0_101));
   AOI21_X1 i_0_0_143 (.A(n_0_0_103), .B1(n_0_0_105), .B2(n_0_0_150), .ZN(
      n_0_0_102));
   INV_X1 i_0_0_144 (.A(n_0_0_104), .ZN(n_0_0_103));
   AOI22_X1 i_0_0_145 (.A1(A[18]), .A2(n_0_0_122), .B1(n_0_0_121), .B2(A[19]), 
      .ZN(n_0_0_104));
   MUX2_X1 i_0_0_146 (.A(A[17]), .B(A[16]), .S(n_0_0_316), .Z(n_0_0_105));
   OAI21_X1 i_0_0_147 (.A(n_0_0_106), .B1(n_0_0_107), .B2(n_0_0_140), .ZN(n_0_66));
   NAND2_X1 i_0_0_148 (.A1(A[17]), .A2(n_0_0_474), .ZN(n_0_0_106));
   MUX2_X1 i_0_0_149 (.A(n_0_0_130), .B(n_0_0_108), .S(n_0_0_146), .Z(n_0_0_107));
   AOI21_X1 i_0_0_150 (.A(n_0_0_109), .B1(n_0_0_111), .B2(n_0_0_150), .ZN(
      n_0_0_108));
   INV_X1 i_0_0_151 (.A(n_0_0_110), .ZN(n_0_0_109));
   AOI22_X1 i_0_0_152 (.A1(A[19]), .A2(n_0_0_122), .B1(n_0_0_121), .B2(A[20]), 
      .ZN(n_0_0_110));
   MUX2_X1 i_0_0_153 (.A(A[18]), .B(A[17]), .S(n_0_0_316), .Z(n_0_0_111));
   OAI21_X1 i_0_0_154 (.A(n_0_0_112), .B1(n_0_0_113), .B2(n_0_0_140), .ZN(n_0_67));
   NAND2_X1 i_0_0_155 (.A1(A[18]), .A2(n_0_0_474), .ZN(n_0_0_112));
   MUX2_X1 i_0_0_156 (.A(n_0_0_135), .B(n_0_0_114), .S(n_0_0_146), .Z(n_0_0_113));
   AOI221_X1 i_0_0_157 (.A(n_0_0_115), .B1(n_0_0_122), .B2(A[20]), .C1(A[21]), 
      .C2(n_0_0_121), .ZN(n_0_0_114));
   INV_X1 i_0_0_158 (.A(n_0_0_116), .ZN(n_0_0_115));
   AOI22_X1 i_0_0_159 (.A1(A[18]), .A2(n_0_0_521), .B1(n_0_0_136), .B2(A[19]), 
      .ZN(n_0_0_116));
   OAI21_X1 i_0_0_160 (.A(n_0_0_117), .B1(n_0_0_118), .B2(n_0_0_140), .ZN(n_0_68));
   NAND2_X1 i_0_0_161 (.A1(A[19]), .A2(n_0_0_474), .ZN(n_0_0_117));
   OAI21_X1 i_0_0_162 (.A(n_0_0_119), .B1(n_0_0_146), .B2(n_0_0_521), .ZN(
      n_0_0_118));
   NAND2_X1 i_0_0_163 (.A1(n_0_0_120), .A2(n_0_0_146), .ZN(n_0_0_119));
   AOI221_X1 i_0_0_164 (.A(n_0_0_124), .B1(n_0_0_122), .B2(A[21]), .C1(n_0_0_121), 
      .C2(A[22]), .ZN(n_0_0_120));
   AND2_X1 i_0_0_165 (.A1(n_0_0_123), .A2(n_0_0_315), .ZN(n_0_0_121));
   AND2_X1 i_0_0_166 (.A1(n_0_0_316), .A2(n_0_0_123), .ZN(n_0_0_122));
   AND2_X1 i_0_0_167 (.A1(n_0_0_152), .A2(n_0_0_151), .ZN(n_0_0_123));
   INV_X1 i_0_0_168 (.A(n_0_0_125), .ZN(n_0_0_124));
   AOI22_X1 i_0_0_169 (.A1(A[19]), .A2(n_0_0_521), .B1(n_0_0_136), .B2(A[20]), 
      .ZN(n_0_0_125));
   OAI21_X1 i_0_0_170 (.A(n_0_0_126), .B1(n_0_0_127), .B2(n_0_0_138), .ZN(n_0_69));
   NAND2_X1 i_0_0_171 (.A1(A[20]), .A2(n_0_0_474), .ZN(n_0_0_126));
   AOI22_X1 i_0_0_172 (.A1(A[20]), .A2(n_0_0_521), .B1(n_0_0_128), .B2(n_0_0_152), 
      .ZN(n_0_0_127));
   OAI21_X1 i_0_0_173 (.A(n_0_0_129), .B1(n_0_0_316), .B2(n_0_0_499), .ZN(
      n_0_0_128));
   OAI21_X1 i_0_0_174 (.A(n_0_0_151), .B1(n_0_0_315), .B2(A[22]), .ZN(n_0_0_129));
   OAI22_X1 i_0_0_175 (.A1(n_0_0_499), .A2(n_0_96), .B1(n_0_0_138), .B2(
      n_0_0_130), .ZN(n_0_70));
   OAI211_X1 i_0_0_176 (.A(n_0_0_152), .B(n_0_0_131), .C1(A[22]), .C2(n_0_0_316), 
      .ZN(n_0_0_130));
   INV_X1 i_0_0_177 (.A(n_0_0_132), .ZN(n_0_0_131));
   MUX2_X1 i_0_0_178 (.A(n_0_0_133), .B(n_0_0_317), .S(n_0_0_314), .Z(n_0_0_132));
   OAI21_X1 i_0_0_179 (.A(n_0_0_497), .B1(n_0_0_317), .B2(A[21]), .ZN(n_0_0_133));
   OAI21_X1 i_0_0_180 (.A(n_0_0_134), .B1(n_0_0_138), .B2(n_0_0_135), .ZN(n_0_71));
   NAND2_X1 i_0_0_181 (.A1(A[22]), .A2(n_0_0_474), .ZN(n_0_0_134));
   OAI21_X1 i_0_0_182 (.A(n_0_0_150), .B1(n_0_0_315), .B2(A[22]), .ZN(n_0_0_135));
   AND2_X1 i_0_0_183 (.A1(n_0_0_150), .A2(n_0_0_315), .ZN(n_0_0_136));
   INV_X1 i_0_0_184 (.A(n_0_0_138), .ZN(n_0_0_137));
   NAND2_X1 i_0_0_185 (.A1(n_0_0_144), .A2(n_0_0_141), .ZN(n_0_0_138));
   INV_X1 i_0_0_186 (.A(n_0_0_140), .ZN(n_0_0_139));
   NAND2_X1 i_0_0_187 (.A1(n_0_0_147), .A2(n_0_0_141), .ZN(n_0_0_140));
   NOR2_X1 i_0_0_188 (.A1(n_0_0_474), .A2(n_0_0_156), .ZN(n_0_0_141));
   OAI21_X1 i_0_0_189 (.A(n_0_96), .B1(n_0_0_156), .B2(n_0_0_142), .ZN(n_0_72));
   NAND2_X1 i_0_0_190 (.A1(n_0_0_521), .A2(n_0_0_144), .ZN(n_0_0_142));
   NAND2_X1 i_0_0_191 (.A1(n_0_0_147), .A2(n_0_0_146), .ZN(n_0_0_143));
   NOR2_X1 i_0_0_192 (.A1(n_0_0_148), .A2(n_0_0_145), .ZN(n_0_0_144));
   INV_X1 i_0_0_193 (.A(n_0_0_146), .ZN(n_0_0_145));
   XNOR2_X1 i_0_0_194 (.A(n_0_0_493), .B(n_0_0_311), .ZN(n_0_0_146));
   INV_X1 i_0_0_195 (.A(n_0_0_148), .ZN(n_0_0_147));
   XNOR2_X1 i_0_0_196 (.A(n_0_0_491), .B(n_0_0_292), .ZN(n_0_0_148));
   NAND2_X1 i_0_0_197 (.A1(n_0_0_316), .A2(n_0_0_150), .ZN(n_0_0_149));
   AOI211_X1 i_0_0_198 (.A(n_0_0_155), .B(n_0_0_151), .C1(n_0_0_153), .C2(
      n_0_0_484), .ZN(n_0_0_150));
   XNOR2_X1 i_0_0_199 (.A(n_0_0_497), .B(n_0_0_314), .ZN(n_0_0_151));
   AOI21_X1 i_0_0_200 (.A(n_0_0_155), .B1(n_0_0_153), .B2(n_0_0_484), .ZN(
      n_0_0_152));
   AOI22_X1 i_0_0_201 (.A1(n_0_0_154), .A2(n_0_0_479), .B1(n_0_0_519), .B2(
      n_0_0_303), .ZN(n_0_0_153));
   MUX2_X1 i_0_0_202 (.A(n_0_0_483), .B(n_0_0_481), .S(n_0_0_309), .Z(n_0_0_154));
   AOI21_X1 i_0_0_203 (.A(n_0_0_484), .B1(n_0_0_303), .B2(n_0_0_300), .ZN(
      n_0_0_155));
   XOR2_X1 i_0_0_204 (.A(n_0_0_487), .B(n_0_0_294), .Z(n_0_0_156));
   OAI221_X1 i_0_0_205 (.A(n_0_0_157), .B1(n_0_0_196), .B2(n_0_0_253), .C1(
      n_0_0_288), .C2(n_0_0_159), .ZN(n_0_73));
   AOI21_X1 i_0_0_206 (.A(n_0_0_158), .B1(n_0_96), .B2(B[0]), .ZN(n_0_0_157));
   NOR2_X1 i_0_0_207 (.A1(n_0_0_246), .A2(n_0_0_211), .ZN(n_0_0_158));
   OAI21_X1 i_0_0_208 (.A(n_0_0_160), .B1(n_0_0_184), .B2(n_0_0_522), .ZN(
      n_0_0_159));
   OAI21_X1 i_0_0_209 (.A(n_0_0_161), .B1(n_0_0_162), .B2(n_0_0_297), .ZN(
      n_0_0_160));
   AOI21_X1 i_0_0_210 (.A(n_0_0_268), .B1(n_0_0_274), .B2(B[3]), .ZN(n_0_0_161));
   AOI22_X1 i_0_0_211 (.A1(n_0_0_163), .A2(n_0_0_316), .B1(B[1]), .B2(n_0_0_281), 
      .ZN(n_0_0_162));
   MUX2_X1 i_0_0_212 (.A(B[2]), .B(B[0]), .S(n_0_0_313), .Z(n_0_0_163));
   OAI21_X1 i_0_0_213 (.A(n_0_0_164), .B1(n_0_0_196), .B2(n_0_0_258), .ZN(n_0_74));
   AOI211_X1 i_0_0_214 (.A(n_0_0_166), .B(n_0_0_165), .C1(B[1]), .C2(n_0_96), 
      .ZN(n_0_0_164));
   NOR2_X1 i_0_0_215 (.A1(n_0_0_246), .A2(n_0_0_216), .ZN(n_0_0_165));
   AOI211_X1 i_0_0_216 (.A(n_0_0_288), .B(n_0_0_167), .C1(n_0_0_191), .C2(
      n_0_0_310), .ZN(n_0_0_166));
   AND3_X1 i_0_0_217 (.A1(n_0_0_169), .A2(n_0_0_168), .A3(n_0_0_522), .ZN(
      n_0_0_167));
   AOI22_X1 i_0_0_218 (.A1(B[4]), .A2(n_0_0_274), .B1(n_0_0_271), .B2(B[3]), 
      .ZN(n_0_0_168));
   AOI22_X1 i_0_0_219 (.A1(B[1]), .A2(n_0_0_275), .B1(n_0_0_273), .B2(B[2]), 
      .ZN(n_0_0_169));
   MUX2_X1 i_0_0_220 (.A(B[2]), .B(n_0_0_170), .S(n_0_0_474), .Z(n_0_75));
   OAI221_X1 i_0_0_221 (.A(n_0_0_171), .B1(n_0_0_210), .B2(n_0_0_262), .C1(
      n_0_0_221), .C2(n_0_0_247), .ZN(n_0_0_170));
   AOI21_X1 i_0_0_222 (.A(n_0_0_172), .B1(n_0_0_199), .B2(n_0_0_204), .ZN(
      n_0_0_171));
   AOI21_X1 i_0_0_223 (.A(n_0_0_206), .B1(n_0_0_174), .B2(n_0_0_173), .ZN(
      n_0_0_172));
   AOI22_X1 i_0_0_224 (.A1(B[2]), .A2(n_0_0_287), .B1(n_0_0_285), .B2(B[5]), 
      .ZN(n_0_0_173));
   AOI22_X1 i_0_0_225 (.A1(B[3]), .A2(n_0_0_281), .B1(n_0_0_279), .B2(B[4]), 
      .ZN(n_0_0_174));
   MUX2_X1 i_0_0_226 (.A(B[3]), .B(n_0_0_175), .S(n_0_0_474), .Z(n_0_76));
   OAI221_X1 i_0_0_227 (.A(n_0_0_176), .B1(n_0_0_226), .B2(n_0_0_247), .C1(
      n_0_0_267), .C2(n_0_0_210), .ZN(n_0_0_175));
   AOI21_X1 i_0_0_228 (.A(n_0_0_177), .B1(n_0_0_204), .B2(n_0_0_207), .ZN(
      n_0_0_176));
   AOI21_X1 i_0_0_229 (.A(n_0_0_206), .B1(n_0_0_179), .B2(n_0_0_178), .ZN(
      n_0_0_177));
   AOI22_X1 i_0_0_230 (.A1(B[3]), .A2(n_0_0_287), .B1(n_0_0_285), .B2(B[6]), 
      .ZN(n_0_0_178));
   AOI22_X1 i_0_0_231 (.A1(B[4]), .A2(n_0_0_281), .B1(n_0_0_279), .B2(B[5]), 
      .ZN(n_0_0_179));
   OAI221_X1 i_0_0_232 (.A(n_0_0_180), .B1(n_0_0_231), .B2(n_0_0_246), .C1(
      n_0_0_288), .C2(n_0_0_182), .ZN(n_0_77));
   AOI21_X1 i_0_0_233 (.A(n_0_0_181), .B1(n_0_96), .B2(B[4]), .ZN(n_0_0_180));
   NOR2_X1 i_0_0_234 (.A1(n_0_0_276), .A2(n_0_0_196), .ZN(n_0_0_181));
   AOI21_X1 i_0_0_235 (.A(n_0_0_183), .B1(n_0_0_184), .B2(n_0_0_522), .ZN(
      n_0_0_182));
   AOI211_X1 i_0_0_236 (.A(n_0_0_522), .B(n_0_0_297), .C1(n_0_0_214), .C2(
      n_0_0_213), .ZN(n_0_0_183));
   NAND2_X1 i_0_0_237 (.A1(n_0_0_186), .A2(n_0_0_185), .ZN(n_0_0_184));
   AOI22_X1 i_0_0_238 (.A1(B[7]), .A2(n_0_0_274), .B1(n_0_0_271), .B2(B[6]), 
      .ZN(n_0_0_185));
   AOI22_X1 i_0_0_239 (.A1(B[4]), .A2(n_0_0_275), .B1(n_0_0_273), .B2(B[5]), 
      .ZN(n_0_0_186));
   OR3_X1 i_0_0_240 (.A1(n_0_0_190), .A2(n_0_0_189), .A3(n_0_0_187), .ZN(n_0_78));
   OAI221_X1 i_0_0_241 (.A(n_0_0_188), .B1(n_0_0_196), .B2(n_0_0_282), .C1(
      n_0_0_236), .C2(n_0_0_246), .ZN(n_0_0_187));
   NAND2_X1 i_0_0_242 (.A1(n_0_96), .A2(B[5]), .ZN(n_0_0_188));
   AND4_X1 i_0_0_243 (.A1(n_0_0_474), .A2(n_0_0_289), .A3(n_0_0_268), .A4(
      n_0_0_217), .ZN(n_0_0_189));
   NOR3_X1 i_0_0_244 (.A1(n_0_0_310), .A2(n_0_0_191), .A3(n_0_0_288), .ZN(
      n_0_0_190));
   AOI221_X1 i_0_0_245 (.A(n_0_0_192), .B1(n_0_0_271), .B2(B[7]), .C1(B[8]), 
      .C2(n_0_0_274), .ZN(n_0_0_191));
   INV_X1 i_0_0_246 (.A(n_0_0_193), .ZN(n_0_0_192));
   AOI22_X1 i_0_0_247 (.A1(B[5]), .A2(n_0_0_275), .B1(n_0_0_273), .B2(B[6]), 
      .ZN(n_0_0_193));
   OAI21_X1 i_0_0_248 (.A(n_0_0_194), .B1(n_0_0_241), .B2(n_0_0_246), .ZN(n_0_79));
   AOI211_X1 i_0_0_249 (.A(n_0_0_197), .B(n_0_0_195), .C1(B[6]), .C2(n_0_96), 
      .ZN(n_0_0_194));
   NOR2_X1 i_0_0_250 (.A1(n_0_0_295), .A2(n_0_0_196), .ZN(n_0_0_195));
   OR2_X1 i_0_0_251 (.A1(n_0_96), .A2(n_0_0_210), .ZN(n_0_0_196));
   NOR2_X1 i_0_0_252 (.A1(n_0_0_288), .A2(n_0_0_198), .ZN(n_0_0_197));
   AOI22_X1 i_0_0_253 (.A1(n_0_0_268), .A2(n_0_0_222), .B1(n_0_0_199), .B2(
      n_0_0_296), .ZN(n_0_0_198));
   NAND2_X1 i_0_0_254 (.A1(n_0_0_201), .A2(n_0_0_200), .ZN(n_0_0_199));
   AOI22_X1 i_0_0_255 (.A1(B[9]), .A2(n_0_0_285), .B1(n_0_0_279), .B2(B[8]), 
      .ZN(n_0_0_200));
   AOI22_X1 i_0_0_256 (.A1(B[6]), .A2(n_0_0_287), .B1(n_0_0_281), .B2(B[7]), 
      .ZN(n_0_0_201));
   MUX2_X1 i_0_0_257 (.A(B[7]), .B(n_0_0_202), .S(n_0_0_474), .Z(n_0_80));
   OAI221_X1 i_0_0_258 (.A(n_0_0_203), .B1(n_0_0_210), .B2(n_0_0_248), .C1(
      n_0_0_249), .C2(n_0_0_247), .ZN(n_0_0_202));
   AOI22_X1 i_0_0_259 (.A1(n_0_0_207), .A2(n_0_0_205), .B1(n_0_0_204), .B2(
      n_0_0_227), .ZN(n_0_0_203));
   AND2_X1 i_0_0_260 (.A1(n_0_0_289), .A2(n_0_0_268), .ZN(n_0_0_204));
   INV_X1 i_0_0_261 (.A(n_0_0_206), .ZN(n_0_0_205));
   NAND2_X1 i_0_0_262 (.A1(n_0_0_296), .A2(n_0_0_289), .ZN(n_0_0_206));
   NAND2_X1 i_0_0_263 (.A1(n_0_0_209), .A2(n_0_0_208), .ZN(n_0_0_207));
   AOI22_X1 i_0_0_264 (.A1(B[10]), .A2(n_0_0_285), .B1(n_0_0_279), .B2(B[9]), 
      .ZN(n_0_0_208));
   AOI22_X1 i_0_0_265 (.A1(B[7]), .A2(n_0_0_287), .B1(n_0_0_281), .B2(B[8]), 
      .ZN(n_0_0_209));
   OR2_X1 i_0_0_266 (.A1(n_0_0_293), .A2(n_0_0_291), .ZN(n_0_0_210));
   OAI221_X1 i_0_0_267 (.A(n_0_0_215), .B1(n_0_0_211), .B2(n_0_0_288), .C1(
      n_0_0_253), .C2(n_0_0_246), .ZN(n_0_81));
   AOI22_X1 i_0_0_268 (.A1(n_0_0_268), .A2(n_0_0_232), .B1(n_0_0_212), .B2(
      n_0_0_296), .ZN(n_0_0_211));
   NAND2_X1 i_0_0_269 (.A1(n_0_0_214), .A2(n_0_0_213), .ZN(n_0_0_212));
   AOI22_X1 i_0_0_270 (.A1(B[11]), .A2(n_0_0_285), .B1(n_0_0_279), .B2(B[10]), 
      .ZN(n_0_0_213));
   AOI22_X1 i_0_0_271 (.A1(B[8]), .A2(n_0_0_287), .B1(n_0_0_281), .B2(B[9]), 
      .ZN(n_0_0_214));
   NAND2_X1 i_0_0_272 (.A1(n_0_96), .A2(B[8]), .ZN(n_0_0_215));
   OAI221_X1 i_0_0_273 (.A(n_0_0_220), .B1(n_0_0_216), .B2(n_0_0_288), .C1(
      n_0_0_258), .C2(n_0_0_246), .ZN(n_0_82));
   AOI22_X1 i_0_0_274 (.A1(n_0_0_296), .A2(n_0_0_217), .B1(n_0_0_268), .B2(
      n_0_0_237), .ZN(n_0_0_216));
   NAND2_X1 i_0_0_275 (.A1(n_0_0_219), .A2(n_0_0_218), .ZN(n_0_0_217));
   AOI22_X1 i_0_0_276 (.A1(B[12]), .A2(n_0_0_285), .B1(n_0_0_279), .B2(B[11]), 
      .ZN(n_0_0_218));
   AOI22_X1 i_0_0_277 (.A1(B[9]), .A2(n_0_0_287), .B1(n_0_0_281), .B2(B[10]), 
      .ZN(n_0_0_219));
   NAND2_X1 i_0_0_278 (.A1(n_0_96), .A2(B[9]), .ZN(n_0_0_220));
   OAI221_X1 i_0_0_279 (.A(n_0_0_225), .B1(n_0_0_246), .B2(n_0_0_262), .C1(
      n_0_0_221), .C2(n_0_0_288), .ZN(n_0_83));
   AOI22_X1 i_0_0_280 (.A1(n_0_0_242), .A2(n_0_0_310), .B1(n_0_0_296), .B2(
      n_0_0_222), .ZN(n_0_0_221));
   NAND2_X1 i_0_0_281 (.A1(n_0_0_224), .A2(n_0_0_223), .ZN(n_0_0_222));
   AOI22_X1 i_0_0_282 (.A1(B[13]), .A2(n_0_0_285), .B1(n_0_0_279), .B2(B[12]), 
      .ZN(n_0_0_223));
   AOI22_X1 i_0_0_283 (.A1(B[10]), .A2(n_0_0_287), .B1(n_0_0_281), .B2(B[11]), 
      .ZN(n_0_0_224));
   NAND2_X1 i_0_0_284 (.A1(n_0_96), .A2(B[10]), .ZN(n_0_0_225));
   OAI221_X1 i_0_0_285 (.A(n_0_0_230), .B1(n_0_0_226), .B2(n_0_0_288), .C1(
      n_0_0_267), .C2(n_0_0_246), .ZN(n_0_84));
   AOI22_X1 i_0_0_286 (.A1(n_0_0_268), .A2(n_0_0_250), .B1(n_0_0_227), .B2(
      n_0_0_296), .ZN(n_0_0_226));
   NAND2_X1 i_0_0_287 (.A1(n_0_0_229), .A2(n_0_0_228), .ZN(n_0_0_227));
   AOI22_X1 i_0_0_288 (.A1(B[14]), .A2(n_0_0_285), .B1(n_0_0_279), .B2(B[13]), 
      .ZN(n_0_0_228));
   AOI22_X1 i_0_0_289 (.A1(B[11]), .A2(n_0_0_287), .B1(n_0_0_281), .B2(B[12]), 
      .ZN(n_0_0_229));
   NAND2_X1 i_0_0_290 (.A1(n_0_96), .A2(B[11]), .ZN(n_0_0_230));
   OAI221_X1 i_0_0_291 (.A(n_0_0_235), .B1(n_0_0_246), .B2(n_0_0_276), .C1(
      n_0_0_231), .C2(n_0_0_288), .ZN(n_0_85));
   AOI22_X1 i_0_0_292 (.A1(n_0_0_254), .A2(n_0_0_310), .B1(n_0_0_296), .B2(
      n_0_0_232), .ZN(n_0_0_231));
   NAND2_X1 i_0_0_293 (.A1(n_0_0_234), .A2(n_0_0_233), .ZN(n_0_0_232));
   AOI22_X1 i_0_0_294 (.A1(B[15]), .A2(n_0_0_285), .B1(n_0_0_279), .B2(B[14]), 
      .ZN(n_0_0_233));
   AOI22_X1 i_0_0_295 (.A1(B[12]), .A2(n_0_0_287), .B1(n_0_0_281), .B2(B[13]), 
      .ZN(n_0_0_234));
   NAND2_X1 i_0_0_296 (.A1(n_0_96), .A2(B[12]), .ZN(n_0_0_235));
   OAI221_X1 i_0_0_297 (.A(n_0_0_240), .B1(n_0_0_246), .B2(n_0_0_282), .C1(
      n_0_0_236), .C2(n_0_0_288), .ZN(n_0_86));
   AOI22_X1 i_0_0_298 (.A1(n_0_0_310), .A2(n_0_0_259), .B1(n_0_0_237), .B2(
      n_0_0_296), .ZN(n_0_0_236));
   NAND2_X1 i_0_0_299 (.A1(n_0_0_239), .A2(n_0_0_238), .ZN(n_0_0_237));
   AOI22_X1 i_0_0_300 (.A1(B[16]), .A2(n_0_0_285), .B1(n_0_0_279), .B2(B[15]), 
      .ZN(n_0_0_238));
   AOI22_X1 i_0_0_301 (.A1(B[13]), .A2(n_0_0_287), .B1(n_0_0_281), .B2(B[14]), 
      .ZN(n_0_0_239));
   NAND2_X1 i_0_0_302 (.A1(n_0_96), .A2(B[13]), .ZN(n_0_0_240));
   OAI221_X1 i_0_0_303 (.A(n_0_0_245), .B1(n_0_0_241), .B2(n_0_0_288), .C1(
      n_0_0_246), .C2(n_0_0_295), .ZN(n_0_87));
   AOI22_X1 i_0_0_304 (.A1(n_0_0_522), .A2(n_0_0_242), .B1(n_0_0_265), .B2(
      n_0_0_268), .ZN(n_0_0_241));
   NAND2_X1 i_0_0_305 (.A1(n_0_0_244), .A2(n_0_0_243), .ZN(n_0_0_242));
   AOI22_X1 i_0_0_306 (.A1(B[17]), .A2(n_0_0_274), .B1(n_0_0_271), .B2(B[16]), 
      .ZN(n_0_0_243));
   AOI22_X1 i_0_0_307 (.A1(B[14]), .A2(n_0_0_275), .B1(n_0_0_273), .B2(B[15]), 
      .ZN(n_0_0_244));
   NAND2_X1 i_0_0_308 (.A1(n_0_96), .A2(B[14]), .ZN(n_0_0_245));
   OAI221_X1 i_0_0_309 (.A(n_0_0_252), .B1(n_0_0_248), .B2(n_0_0_246), .C1(
      n_0_0_249), .C2(n_0_0_288), .ZN(n_0_88));
   OR2_X1 i_0_0_310 (.A1(n_0_96), .A2(n_0_0_247), .ZN(n_0_0_246));
   NAND2_X1 i_0_0_311 (.A1(n_0_0_293), .A2(n_0_0_291), .ZN(n_0_0_247));
   NAND2_X1 i_0_0_312 (.A1(n_0_0_296), .A2(n_0_0_287), .ZN(n_0_0_248));
   AOI22_X1 i_0_0_313 (.A1(n_0_0_269), .A2(n_0_0_310), .B1(n_0_0_296), .B2(
      n_0_0_250), .ZN(n_0_0_249));
   OAI221_X1 i_0_0_314 (.A(n_0_0_251), .B1(n_0_0_278), .B2(n_0_0_505), .C1(
      n_0_0_506), .C2(n_0_0_284), .ZN(n_0_0_250));
   AOI22_X1 i_0_0_315 (.A1(B[15]), .A2(n_0_0_287), .B1(n_0_0_281), .B2(B[16]), 
      .ZN(n_0_0_251));
   NAND2_X1 i_0_0_316 (.A1(n_0_96), .A2(B[15]), .ZN(n_0_0_252));
   OAI21_X1 i_0_0_317 (.A(n_0_0_257), .B1(n_0_0_253), .B2(n_0_0_288), .ZN(n_0_89));
   AOI22_X1 i_0_0_318 (.A1(n_0_0_522), .A2(n_0_0_254), .B1(n_0_0_268), .B2(
      n_0_0_277), .ZN(n_0_0_253));
   NAND2_X1 i_0_0_319 (.A1(n_0_0_256), .A2(n_0_0_255), .ZN(n_0_0_254));
   AOI22_X1 i_0_0_320 (.A1(B[19]), .A2(n_0_0_274), .B1(n_0_0_271), .B2(B[18]), 
      .ZN(n_0_0_255));
   AOI22_X1 i_0_0_321 (.A1(B[16]), .A2(n_0_0_275), .B1(n_0_0_273), .B2(B[17]), 
      .ZN(n_0_0_256));
   NAND2_X1 i_0_0_322 (.A1(n_0_96), .A2(B[16]), .ZN(n_0_0_257));
   OAI22_X1 i_0_0_323 (.A1(n_0_0_288), .A2(n_0_0_258), .B1(n_0_0_505), .B2(
      n_0_0_474), .ZN(n_0_90));
   AOI22_X1 i_0_0_324 (.A1(n_0_0_522), .A2(n_0_0_259), .B1(n_0_0_268), .B2(
      n_0_0_283), .ZN(n_0_0_258));
   NAND2_X1 i_0_0_325 (.A1(n_0_0_261), .A2(n_0_0_260), .ZN(n_0_0_259));
   AOI22_X1 i_0_0_326 (.A1(B[20]), .A2(n_0_0_274), .B1(n_0_0_271), .B2(B[19]), 
      .ZN(n_0_0_260));
   AOI22_X1 i_0_0_327 (.A1(B[17]), .A2(n_0_0_275), .B1(n_0_0_273), .B2(B[18]), 
      .ZN(n_0_0_261));
   OAI22_X1 i_0_0_328 (.A1(n_0_0_288), .A2(n_0_0_262), .B1(n_0_0_506), .B2(
      n_0_0_474), .ZN(n_0_91));
   AOI21_X1 i_0_0_329 (.A(n_0_0_263), .B1(n_0_0_265), .B2(n_0_0_296), .ZN(
      n_0_0_262));
   NOR3_X1 i_0_0_330 (.A1(n_0_0_523), .A2(n_0_0_297), .A3(n_0_0_264), .ZN(
      n_0_0_263));
   OAI21_X1 i_0_0_331 (.A(n_0_0_310), .B1(n_0_0_315), .B2(B[22]), .ZN(n_0_0_264));
   OAI221_X1 i_0_0_332 (.A(n_0_0_266), .B1(n_0_0_286), .B2(n_0_0_506), .C1(
      n_0_0_507), .C2(n_0_0_280), .ZN(n_0_0_265));
   AOI22_X1 i_0_0_333 (.A1(B[21]), .A2(n_0_0_285), .B1(n_0_0_279), .B2(B[20]), 
      .ZN(n_0_0_266));
   OAI22_X1 i_0_0_334 (.A1(n_0_0_288), .A2(n_0_0_267), .B1(n_0_0_507), .B2(
      n_0_0_474), .ZN(n_0_92));
   AOI22_X1 i_0_0_335 (.A1(n_0_0_522), .A2(n_0_0_269), .B1(n_0_0_268), .B2(
      n_0_0_287), .ZN(n_0_0_267));
   NOR2_X1 i_0_0_336 (.A1(n_0_0_297), .A2(n_0_0_522), .ZN(n_0_0_268));
   NAND2_X1 i_0_0_337 (.A1(n_0_0_272), .A2(n_0_0_270), .ZN(n_0_0_269));
   AOI22_X1 i_0_0_338 (.A1(B[22]), .A2(n_0_0_274), .B1(n_0_0_271), .B2(B[21]), 
      .ZN(n_0_0_270));
   NOR2_X1 i_0_0_339 (.A1(n_0_0_297), .A2(n_0_0_278), .ZN(n_0_0_271));
   AOI22_X1 i_0_0_340 (.A1(B[19]), .A2(n_0_0_275), .B1(n_0_0_273), .B2(B[20]), 
      .ZN(n_0_0_272));
   NOR2_X1 i_0_0_341 (.A1(n_0_0_297), .A2(n_0_0_280), .ZN(n_0_0_273));
   NOR2_X1 i_0_0_342 (.A1(n_0_0_297), .A2(n_0_0_284), .ZN(n_0_0_274));
   NOR2_X1 i_0_0_343 (.A1(n_0_0_297), .A2(n_0_0_286), .ZN(n_0_0_275));
   OAI22_X1 i_0_0_344 (.A1(n_0_0_288), .A2(n_0_0_276), .B1(n_0_0_508), .B2(
      n_0_0_474), .ZN(n_0_93));
   NAND2_X1 i_0_0_345 (.A1(n_0_0_296), .A2(n_0_0_277), .ZN(n_0_0_276));
   AOI222_X1 i_0_0_346 (.A1(n_0_0_281), .A2(n_0_0_509), .B1(n_0_0_287), .B2(
      n_0_0_508), .C1(n_0_0_279), .C2(n_0_0_510), .ZN(n_0_0_277));
   NAND2_X1 i_0_0_347 (.A1(n_0_0_316), .A2(n_0_0_523), .ZN(n_0_0_278));
   NOR2_X1 i_0_0_348 (.A1(n_0_0_315), .A2(n_0_0_313), .ZN(n_0_0_279));
   NAND2_X1 i_0_0_349 (.A1(n_0_0_315), .A2(n_0_0_313), .ZN(n_0_0_280));
   NOR2_X1 i_0_0_350 (.A1(n_0_0_316), .A2(n_0_0_523), .ZN(n_0_0_281));
   OAI22_X1 i_0_0_351 (.A1(n_0_0_288), .A2(n_0_0_282), .B1(n_0_0_509), .B2(
      n_0_0_474), .ZN(n_0_94));
   NAND2_X1 i_0_0_352 (.A1(n_0_0_296), .A2(n_0_0_283), .ZN(n_0_0_282));
   AOI221_X1 i_0_0_353 (.A(n_0_0_285), .B1(n_0_0_315), .B2(n_0_0_510), .C1(
      n_0_0_287), .C2(n_0_0_509), .ZN(n_0_0_283));
   INV_X1 i_0_0_354 (.A(n_0_0_285), .ZN(n_0_0_284));
   NOR2_X1 i_0_0_355 (.A1(n_0_0_313), .A2(n_0_0_316), .ZN(n_0_0_285));
   INV_X1 i_0_0_356 (.A(n_0_0_287), .ZN(n_0_0_286));
   NOR2_X1 i_0_0_357 (.A1(n_0_0_523), .A2(n_0_0_315), .ZN(n_0_0_287));
   OAI22_X1 i_0_0_358 (.A1(n_0_0_295), .A2(n_0_0_288), .B1(n_0_0_510), .B2(
      n_0_0_474), .ZN(n_0_95));
   NAND2_X1 i_0_0_359 (.A1(n_0_0_474), .A2(n_0_0_289), .ZN(n_0_0_288));
   AND2_X1 i_0_0_360 (.A1(n_0_0_293), .A2(n_0_0_290), .ZN(n_0_0_289));
   INV_X1 i_0_0_361 (.A(n_0_0_291), .ZN(n_0_0_290));
   XOR2_X1 i_0_0_362 (.A(n_0_0_308), .B(n_0_0_292), .Z(n_0_0_291));
   XNOR2_X1 i_0_0_363 (.A(n_0_0_513), .B(A[26]), .ZN(n_0_0_292));
   XOR2_X1 i_0_0_364 (.A(n_0_0_307), .B(n_0_0_294), .Z(n_0_0_293));
   XNOR2_X1 i_0_0_365 (.A(B[27]), .B(n_0_0_501), .ZN(n_0_0_294));
   OAI211_X1 i_0_0_366 (.A(n_0_0_296), .B(n_0_0_313), .C1(n_0_0_315), .C2(B[22]), 
      .ZN(n_0_0_295));
   NOR2_X1 i_0_0_367 (.A1(n_0_0_310), .A2(n_0_0_297), .ZN(n_0_0_296));
   AOI21_X1 i_0_0_368 (.A(n_0_0_298), .B1(n_0_0_301), .B2(n_0_0_306), .ZN(
      n_0_0_297));
   NOR2_X1 i_0_0_369 (.A1(n_0_0_306), .A2(n_0_0_299), .ZN(n_0_0_298));
   NAND2_X1 i_0_0_370 (.A1(n_0_0_303), .A2(n_0_0_300), .ZN(n_0_0_299));
   NOR2_X1 i_0_0_371 (.A1(n_0_0_519), .A2(n_0_0_479), .ZN(n_0_0_300));
   OAI21_X1 i_0_0_372 (.A(n_0_0_302), .B1(n_0_0_304), .B2(n_0_0_482), .ZN(
      n_0_0_301));
   NAND2_X1 i_0_0_373 (.A1(n_0_0_479), .A2(n_0_0_303), .ZN(n_0_0_302));
   NOR3_X1 i_0_0_374 (.A1(n_0_0_309), .A2(n_0_0_481), .A3(n_0_0_483), .ZN(
      n_0_0_303));
   AOI21_X1 i_0_0_375 (.A(n_0_0_305), .B1(n_0_0_309), .B2(n_0_0_483), .ZN(
      n_0_0_304));
   NOR2_X1 i_0_0_376 (.A1(n_0_0_480), .A2(n_0_0_309), .ZN(n_0_0_305));
   AOI21_X1 i_0_0_377 (.A(n_0_0_490), .B1(n_0_0_307), .B2(n_0_0_486), .ZN(
      n_0_0_306));
   AOI21_X1 i_0_0_378 (.A(n_0_0_488), .B1(n_0_0_308), .B2(n_0_0_489), .ZN(
      n_0_0_307));
   AOI21_X1 i_0_0_379 (.A(n_0_0_495), .B1(n_0_0_492), .B2(n_0_0_312), .ZN(
      n_0_0_308));
   XNOR2_X1 i_0_0_380 (.A(B[30]), .B(n_0_0_504), .ZN(n_0_0_309));
   XNOR2_X1 i_0_0_381 (.A(n_0_0_312), .B(n_0_0_311), .ZN(n_0_0_310));
   XNOR2_X1 i_0_0_382 (.A(B[25]), .B(n_0_0_500), .ZN(n_0_0_311));
   OAI21_X1 i_0_0_383 (.A(n_0_0_496), .B1(n_0_0_494), .B2(n_0_0_317), .ZN(
      n_0_0_312));
   XNOR2_X1 i_0_0_384 (.A(n_0_0_317), .B(n_0_0_314), .ZN(n_0_0_313));
   XNOR2_X1 i_0_0_385 (.A(n_0_0_512), .B(A[24]), .ZN(n_0_0_314));
   XNOR2_X1 i_0_0_386 (.A(n_0_0_511), .B(A[23]), .ZN(n_0_0_315));
   XNOR2_X1 i_0_0_387 (.A(B[23]), .B(A[23]), .ZN(n_0_0_316));
   NOR2_X1 i_0_0_388 (.A1(n_0_0_511), .A2(A[23]), .ZN(n_0_0_317));
   INV_X1 i_0_0_389 (.A(n_0_0_318), .ZN(Sum[0]));
   AOI22_X1 i_0_0_390 (.A1(n_0_1), .A2(n_0_0_527), .B1(n_0_0_526), .B2(n_0_0), 
      .ZN(n_0_0_318));
   OAI21_X1 i_0_0_391 (.A(n_0_0_321), .B1(n_0_0_319), .B2(n_0_0_520), .ZN(Sum[1]));
   AOI21_X1 i_0_0_392 (.A(n_0_0_320), .B1(n_0_2), .B2(n_0_24), .ZN(n_0_0_319));
   NOR2_X1 i_0_0_393 (.A1(n_0_0_515), .A2(n_0_24), .ZN(n_0_0_320));
   NAND3_X1 i_0_0_394 (.A1(n_0_0), .A2(n_0_0_420), .A3(n_0_0_331), .ZN(n_0_0_321));
   OAI21_X1 i_0_0_395 (.A(n_0_0_322), .B1(n_0_0_323), .B2(n_0_0_330), .ZN(Sum[2]));
   AOI22_X1 i_0_0_396 (.A1(n_0_3), .A2(n_0_0_527), .B1(n_0_0_526), .B2(n_0_2), 
      .ZN(n_0_0_322));
   AOI22_X1 i_0_0_397 (.A1(n_0_1), .A2(n_0_0_420), .B1(n_0_0_524), .B2(n_0_0), 
      .ZN(n_0_0_323));
   OAI211_X1 i_0_0_398 (.A(n_0_0_325), .B(n_0_0_324), .C1(n_0_0_525), .C2(
      n_0_0_327), .ZN(Sum[3]));
   AOI22_X1 i_0_0_399 (.A1(n_0_4), .A2(n_0_0_527), .B1(n_0_0_526), .B2(n_0_3), 
      .ZN(n_0_0_324));
   NAND3_X1 i_0_0_400 (.A1(n_0_1), .A2(n_0_0_524), .A3(n_0_0_331), .ZN(n_0_0_325));
   OAI221_X1 i_0_0_401 (.A(n_0_0_326), .B1(n_0_0_327), .B2(n_0_0_419), .C1(
      n_0_0_525), .C2(n_0_0_329), .ZN(Sum[4]));
   AOI22_X1 i_0_0_402 (.A1(n_0_5), .A2(n_0_0_527), .B1(n_0_0_526), .B2(n_0_4), 
      .ZN(n_0_0_326));
   AOI22_X1 i_0_0_403 (.A1(n_0_0), .A2(n_0_0_337), .B1(n_0_0_331), .B2(n_0_2), 
      .ZN(n_0_0_327));
   OAI221_X1 i_0_0_404 (.A(n_0_0_328), .B1(n_0_0_329), .B2(n_0_0_419), .C1(
      n_0_0_525), .C2(n_0_0_332), .ZN(Sum[5]));
   AOI22_X1 i_0_0_405 (.A1(n_0_6), .A2(n_0_0_527), .B1(n_0_0_526), .B2(n_0_5), 
      .ZN(n_0_0_328));
   AOI22_X1 i_0_0_406 (.A1(n_0_1), .A2(n_0_0_337), .B1(n_0_0_331), .B2(n_0_3), 
      .ZN(n_0_0_329));
   INV_X1 i_0_0_407 (.A(n_0_0_331), .ZN(n_0_0_330));
   NOR4_X1 i_0_0_408 (.A1(num_leading_zeros[4]), .A2(num_leading_zeros[3]), 
      .A3(num_leading_zeros[2]), .A4(num_leading_zeros[1]), .ZN(n_0_0_331));
   AOI221_X1 i_0_0_409 (.A(n_0_0_334), .B1(n_0_0_332), .B2(n_0_0_524), .C1(
      n_0_0_335), .C2(n_0_0_420), .ZN(Sum[6]));
   AOI21_X1 i_0_0_410 (.A(n_0_0_333), .B1(n_0_0_337), .B2(n_0_2), .ZN(n_0_0_332));
   NOR2_X1 i_0_0_411 (.A1(n_0_0_340), .A2(num_leading_zeros[1]), .ZN(n_0_0_333));
   OAI22_X1 i_0_0_412 (.A1(n_0_0_387), .A2(n_0_6), .B1(n_0_7), .B2(n_0_0_388), 
      .ZN(n_0_0_334));
   AOI221_X1 i_0_0_413 (.A(n_0_0_338), .B1(n_0_0_335), .B2(n_0_0_524), .C1(
      n_0_0_339), .C2(n_0_0_420), .ZN(Sum[7]));
   AOI21_X1 i_0_0_414 (.A(n_0_0_336), .B1(n_0_0_337), .B2(n_0_3), .ZN(n_0_0_335));
   NOR2_X1 i_0_0_415 (.A1(n_0_0_343), .A2(num_leading_zeros[1]), .ZN(n_0_0_336));
   AND2_X1 i_0_0_416 (.A1(num_leading_zeros[1]), .A2(n_0_0_413), .ZN(n_0_0_337));
   OAI22_X1 i_0_0_417 (.A1(n_0_0_387), .A2(n_0_7), .B1(n_0_8), .B2(n_0_0_388), 
      .ZN(n_0_0_338));
   OAI221_X1 i_0_0_418 (.A(n_0_0_341), .B1(n_0_0_339), .B2(n_0_0_419), .C1(
      n_0_0_342), .C2(n_0_0_525), .ZN(Sum[8]));
   MUX2_X1 i_0_0_419 (.A(n_0_0_346), .B(n_0_0_340), .S(num_leading_zeros[1]), 
      .Z(n_0_0_339));
   AOI22_X1 i_0_0_420 (.A1(n_0_4), .A2(n_0_0_413), .B1(n_0_0_377), .B2(n_0_0), 
      .ZN(n_0_0_340));
   AOI22_X1 i_0_0_421 (.A1(n_0_9), .A2(n_0_0_527), .B1(n_0_0_526), .B2(n_0_8), 
      .ZN(n_0_0_341));
   OAI221_X1 i_0_0_422 (.A(n_0_0_344), .B1(n_0_0_342), .B2(n_0_0_419), .C1(
      n_0_0_345), .C2(n_0_0_525), .ZN(Sum[9]));
   MUX2_X1 i_0_0_423 (.A(n_0_0_349), .B(n_0_0_343), .S(num_leading_zeros[1]), 
      .Z(n_0_0_342));
   AOI22_X1 i_0_0_424 (.A1(n_0_5), .A2(n_0_0_413), .B1(n_0_0_377), .B2(n_0_1), 
      .ZN(n_0_0_343));
   AOI22_X1 i_0_0_425 (.A1(n_0_10), .A2(n_0_0_527), .B1(n_0_0_526), .B2(n_0_9), 
      .ZN(n_0_0_344));
   OAI221_X1 i_0_0_426 (.A(n_0_0_347), .B1(n_0_0_345), .B2(n_0_0_419), .C1(
      n_0_0_348), .C2(n_0_0_525), .ZN(Sum[10]));
   MUX2_X1 i_0_0_427 (.A(n_0_0_352), .B(n_0_0_346), .S(num_leading_zeros[1]), 
      .Z(n_0_0_345));
   AOI22_X1 i_0_0_428 (.A1(n_0_6), .A2(n_0_0_413), .B1(n_0_0_377), .B2(n_0_2), 
      .ZN(n_0_0_346));
   AOI22_X1 i_0_0_429 (.A1(n_0_11), .A2(n_0_0_527), .B1(n_0_0_526), .B2(n_0_10), 
      .ZN(n_0_0_347));
   OAI221_X1 i_0_0_430 (.A(n_0_0_350), .B1(n_0_0_348), .B2(n_0_0_419), .C1(
      n_0_0_351), .C2(n_0_0_525), .ZN(Sum[11]));
   MUX2_X1 i_0_0_431 (.A(n_0_0_355), .B(n_0_0_349), .S(num_leading_zeros[1]), 
      .Z(n_0_0_348));
   AOI22_X1 i_0_0_432 (.A1(n_0_7), .A2(n_0_0_413), .B1(n_0_0_377), .B2(n_0_3), 
      .ZN(n_0_0_349));
   AOI22_X1 i_0_0_433 (.A1(n_0_12), .A2(n_0_0_527), .B1(n_0_0_526), .B2(n_0_11), 
      .ZN(n_0_0_350));
   OAI221_X1 i_0_0_434 (.A(n_0_0_353), .B1(n_0_0_351), .B2(n_0_0_419), .C1(
      n_0_0_354), .C2(n_0_0_525), .ZN(Sum[12]));
   MUX2_X1 i_0_0_435 (.A(n_0_0_359), .B(n_0_0_352), .S(num_leading_zeros[1]), 
      .Z(n_0_0_351));
   AOI222_X1 i_0_0_436 (.A1(n_0_8), .A2(n_0_0_413), .B1(n_0_0_412), .B2(n_0_0), 
      .C1(n_0_0_377), .C2(n_0_4), .ZN(n_0_0_352));
   AOI22_X1 i_0_0_437 (.A1(n_0_13), .A2(n_0_0_527), .B1(n_0_0_526), .B2(n_0_12), 
      .ZN(n_0_0_353));
   OAI221_X1 i_0_0_438 (.A(n_0_0_356), .B1(n_0_0_354), .B2(n_0_0_419), .C1(
      n_0_0_358), .C2(n_0_0_525), .ZN(Sum[13]));
   MUX2_X1 i_0_0_439 (.A(n_0_0_361), .B(n_0_0_355), .S(num_leading_zeros[1]), 
      .Z(n_0_0_354));
   AOI222_X1 i_0_0_440 (.A1(n_0_9), .A2(n_0_0_413), .B1(n_0_0_412), .B2(n_0_1), 
      .C1(n_0_0_377), .C2(n_0_5), .ZN(n_0_0_355));
   AOI22_X1 i_0_0_441 (.A1(n_0_14), .A2(n_0_0_527), .B1(n_0_0_526), .B2(n_0_13), 
      .ZN(n_0_0_356));
   AOI221_X1 i_0_0_442 (.A(n_0_0_357), .B1(n_0_0_358), .B2(n_0_0_524), .C1(
      n_0_0_420), .C2(n_0_0_360), .ZN(Sum[14]));
   OAI22_X1 i_0_0_443 (.A1(n_0_0_387), .A2(n_0_14), .B1(n_0_15), .B2(n_0_0_388), 
      .ZN(n_0_0_357));
   MUX2_X1 i_0_0_444 (.A(n_0_0_365), .B(n_0_0_359), .S(num_leading_zeros[1]), 
      .Z(n_0_0_358));
   AOI222_X1 i_0_0_445 (.A1(n_0_10), .A2(n_0_0_413), .B1(n_0_0_412), .B2(n_0_2), 
      .C1(n_0_0_377), .C2(n_0_6), .ZN(n_0_0_359));
   OAI221_X1 i_0_0_446 (.A(n_0_0_362), .B1(n_0_0_360), .B2(n_0_0_419), .C1(
      n_0_0_364), .C2(n_0_0_525), .ZN(Sum[15]));
   MUX2_X1 i_0_0_447 (.A(n_0_0_369), .B(n_0_0_361), .S(num_leading_zeros[1]), 
      .Z(n_0_0_360));
   AOI222_X1 i_0_0_448 (.A1(n_0_11), .A2(n_0_0_413), .B1(n_0_0_412), .B2(n_0_3), 
      .C1(n_0_0_377), .C2(n_0_7), .ZN(n_0_0_361));
   AOI22_X1 i_0_0_449 (.A1(n_0_16), .A2(n_0_0_527), .B1(n_0_0_526), .B2(n_0_15), 
      .ZN(n_0_0_362));
   OAI221_X1 i_0_0_450 (.A(n_0_0_363), .B1(n_0_0_364), .B2(n_0_0_419), .C1(
      n_0_0_525), .C2(n_0_0_368), .ZN(Sum[16]));
   AOI22_X1 i_0_0_451 (.A1(n_0_17), .A2(n_0_0_527), .B1(n_0_0_526), .B2(n_0_16), 
      .ZN(n_0_0_363));
   MUX2_X1 i_0_0_452 (.A(n_0_0_373), .B(n_0_0_365), .S(num_leading_zeros[1]), 
      .Z(n_0_0_364));
   AOI221_X1 i_0_0_453 (.A(n_0_0_366), .B1(n_0_0_378), .B2(n_0_0), .C1(n_0_8), 
      .C2(n_0_0_377), .ZN(n_0_0_365));
   NOR2_X1 i_0_0_454 (.A1(n_0_0_382), .A2(num_leading_zeros[2]), .ZN(n_0_0_366));
   OAI221_X1 i_0_0_455 (.A(n_0_0_367), .B1(n_0_0_368), .B2(n_0_0_419), .C1(
      n_0_0_525), .C2(n_0_0_372), .ZN(Sum[17]));
   AOI22_X1 i_0_0_456 (.A1(n_0_18), .A2(n_0_0_527), .B1(n_0_0_526), .B2(n_0_17), 
      .ZN(n_0_0_367));
   MUX2_X1 i_0_0_457 (.A(n_0_0_376), .B(n_0_0_369), .S(num_leading_zeros[1]), 
      .Z(n_0_0_368));
   AOI221_X1 i_0_0_458 (.A(n_0_0_370), .B1(n_0_0_378), .B2(n_0_1), .C1(n_0_9), 
      .C2(n_0_0_377), .ZN(n_0_0_369));
   NOR2_X1 i_0_0_459 (.A1(n_0_0_385), .A2(num_leading_zeros[2]), .ZN(n_0_0_370));
   OAI221_X1 i_0_0_460 (.A(n_0_0_371), .B1(n_0_0_372), .B2(n_0_0_419), .C1(
      n_0_0_525), .C2(n_0_0_375), .ZN(Sum[18]));
   AOI22_X1 i_0_0_461 (.A1(n_0_19), .A2(n_0_0_527), .B1(n_0_0_526), .B2(n_0_18), 
      .ZN(n_0_0_371));
   MUX2_X1 i_0_0_462 (.A(n_0_0_381), .B(n_0_0_373), .S(num_leading_zeros[1]), 
      .Z(n_0_0_372));
   AOI222_X1 i_0_0_463 (.A1(n_0_0_414), .A2(n_0_0_516), .B1(n_0_2), .B2(
      n_0_0_378), .C1(n_0_0_377), .C2(n_0_10), .ZN(n_0_0_373));
   OAI221_X1 i_0_0_464 (.A(n_0_0_374), .B1(n_0_0_380), .B2(n_0_0_525), .C1(
      n_0_0_419), .C2(n_0_0_375), .ZN(Sum[19]));
   AOI22_X1 i_0_0_465 (.A1(n_0_20), .A2(n_0_0_527), .B1(n_0_0_526), .B2(n_0_19), 
      .ZN(n_0_0_374));
   MUX2_X1 i_0_0_466 (.A(n_0_0_384), .B(n_0_0_376), .S(num_leading_zeros[1]), 
      .Z(n_0_0_375));
   AOI222_X1 i_0_0_467 (.A1(n_0_0_400), .A2(n_0_0_516), .B1(n_0_3), .B2(
      n_0_0_378), .C1(n_0_0_377), .C2(n_0_11), .ZN(n_0_0_376));
   NOR3_X1 i_0_0_468 (.A1(n_0_0_516), .A2(num_leading_zeros[3]), .A3(
      num_leading_zeros[4]), .ZN(n_0_0_377));
   NOR3_X1 i_0_0_469 (.A1(n_0_0_517), .A2(n_0_0_516), .A3(num_leading_zeros[4]), 
      .ZN(n_0_0_378));
   OAI221_X1 i_0_0_470 (.A(n_0_0_379), .B1(n_0_0_380), .B2(n_0_0_419), .C1(
      n_0_0_525), .C2(n_0_0_383), .ZN(Sum[20]));
   AOI22_X1 i_0_0_471 (.A1(n_0_21), .A2(n_0_0_527), .B1(n_0_0_526), .B2(n_0_20), 
      .ZN(n_0_0_379));
   MUX2_X1 i_0_0_472 (.A(n_0_0_408), .B(n_0_0_381), .S(num_leading_zeros[1]), 
      .Z(n_0_0_380));
   MUX2_X1 i_0_0_473 (.A(n_0_0_382), .B(n_0_0_406), .S(n_0_0_516), .Z(n_0_0_381));
   AOI22_X1 i_0_0_474 (.A1(n_0_4), .A2(n_0_0_417), .B1(n_0_0_416), .B2(n_0_12), 
      .ZN(n_0_0_382));
   AOI221_X1 i_0_0_475 (.A(n_0_0_386), .B1(n_0_0_383), .B2(n_0_0_524), .C1(
      n_0_0_402), .C2(n_0_0_420), .ZN(Sum[21]));
   MUX2_X1 i_0_0_476 (.A(n_0_0_397), .B(n_0_0_384), .S(num_leading_zeros[1]), 
      .Z(n_0_0_383));
   MUX2_X1 i_0_0_477 (.A(n_0_0_385), .B(n_0_0_395), .S(n_0_0_516), .Z(n_0_0_384));
   AOI22_X1 i_0_0_478 (.A1(n_0_5), .A2(n_0_0_417), .B1(n_0_0_416), .B2(n_0_13), 
      .ZN(n_0_0_385));
   OAI22_X1 i_0_0_479 (.A1(n_0_0_387), .A2(n_0_21), .B1(n_0_22), .B2(n_0_0_388), 
      .ZN(n_0_0_386));
   OR2_X1 i_0_0_480 (.A1(n_0_0_520), .A2(n_0_24), .ZN(n_0_0_387));
   NAND2_X1 i_0_0_481 (.A1(n_0_24), .A2(n_0_0_442), .ZN(n_0_0_388));
   AOI21_X1 i_0_0_482 (.A(n_0_0_389), .B1(n_0_0_402), .B2(n_0_0_524), .ZN(
      Sum[22]));
   OAI22_X1 i_0_0_483 (.A1(n_0_0_525), .A2(n_0_0_391), .B1(n_0_0_390), .B2(
      n_0_0_520), .ZN(n_0_0_389));
   MUX2_X1 i_0_0_484 (.A(n_0_22), .B(n_0_23), .S(n_0_24), .Z(n_0_0_390));
   AOI21_X1 i_0_0_485 (.A(n_0_0_392), .B1(n_0_0_397), .B2(num_leading_zeros[1]), 
      .ZN(n_0_0_391));
   NOR2_X1 i_0_0_486 (.A1(num_leading_zeros[1]), .A2(n_0_0_393), .ZN(n_0_0_392));
   OAI21_X1 i_0_0_487 (.A(n_0_0_394), .B1(n_0_0_395), .B2(n_0_0_516), .ZN(
      n_0_0_393));
   AOI222_X1 i_0_0_488 (.A1(n_0_21), .A2(n_0_0_413), .B1(n_0_0_412), .B2(n_0_13), 
      .C1(n_0_0_411), .C2(n_0_5), .ZN(n_0_0_394));
   AOI221_X1 i_0_0_489 (.A(n_0_0_396), .B1(n_0_0_417), .B2(n_0_9), .C1(n_0_17), 
      .C2(n_0_0_416), .ZN(n_0_0_395));
   NOR3_X1 i_0_0_490 (.A1(n_0_0_518), .A2(n_0_0_515), .A3(num_leading_zeros[3]), 
      .ZN(n_0_0_396));
   AOI221_X1 i_0_0_491 (.A(n_0_0_398), .B1(n_0_0_413), .B2(n_0_19), .C1(
      num_leading_zeros[2]), .C2(n_0_0_400), .ZN(n_0_0_397));
   INV_X1 i_0_0_492 (.A(n_0_0_399), .ZN(n_0_0_398));
   AOI22_X1 i_0_0_493 (.A1(n_0_11), .A2(n_0_0_412), .B1(n_0_0_411), .B2(n_0_3), 
      .ZN(n_0_0_399));
   INV_X1 i_0_0_494 (.A(n_0_0_401), .ZN(n_0_0_400));
   AOI22_X1 i_0_0_495 (.A1(n_0_7), .A2(n_0_0_417), .B1(n_0_0_416), .B2(n_0_15), 
      .ZN(n_0_0_401));
   OAI21_X1 i_0_0_496 (.A(n_0_0_403), .B1(n_0_0_404), .B2(num_leading_zeros[1]), 
      .ZN(n_0_0_402));
   NAND2_X1 i_0_0_497 (.A1(n_0_0_408), .A2(num_leading_zeros[1]), .ZN(n_0_0_403));
   OAI21_X1 i_0_0_498 (.A(n_0_0_405), .B1(n_0_0_406), .B2(n_0_0_516), .ZN(
      n_0_0_404));
   AOI222_X1 i_0_0_499 (.A1(n_0_20), .A2(n_0_0_413), .B1(n_0_0_412), .B2(n_0_12), 
      .C1(n_0_0_411), .C2(n_0_4), .ZN(n_0_0_405));
   AOI221_X1 i_0_0_500 (.A(n_0_0_407), .B1(n_0_0_417), .B2(n_0_8), .C1(n_0_16), 
      .C2(n_0_0_416), .ZN(n_0_0_406));
   AND3_X1 i_0_0_501 (.A1(n_0_0_517), .A2(n_0_0), .A3(num_leading_zeros[4]), 
      .ZN(n_0_0_407));
   AOI221_X1 i_0_0_502 (.A(n_0_0_409), .B1(n_0_0_413), .B2(n_0_18), .C1(
      num_leading_zeros[2]), .C2(n_0_0_414), .ZN(n_0_0_408));
   INV_X1 i_0_0_503 (.A(n_0_0_410), .ZN(n_0_0_409));
   AOI22_X1 i_0_0_504 (.A1(n_0_10), .A2(n_0_0_412), .B1(n_0_0_411), .B2(n_0_2), 
      .ZN(n_0_0_410));
   NOR3_X1 i_0_0_505 (.A1(n_0_0_518), .A2(num_leading_zeros[3]), .A3(
      num_leading_zeros[2]), .ZN(n_0_0_411));
   NOR3_X1 i_0_0_506 (.A1(n_0_0_517), .A2(num_leading_zeros[2]), .A3(
      num_leading_zeros[4]), .ZN(n_0_0_412));
   NOR3_X1 i_0_0_507 (.A1(num_leading_zeros[4]), .A2(num_leading_zeros[3]), 
      .A3(num_leading_zeros[2]), .ZN(n_0_0_413));
   INV_X1 i_0_0_508 (.A(n_0_0_415), .ZN(n_0_0_414));
   AOI22_X1 i_0_0_509 (.A1(n_0_6), .A2(n_0_0_417), .B1(n_0_0_416), .B2(n_0_14), 
      .ZN(n_0_0_415));
   NOR2_X1 i_0_0_510 (.A1(num_leading_zeros[4]), .A2(num_leading_zeros[3]), 
      .ZN(n_0_0_416));
   NOR2_X1 i_0_0_511 (.A1(n_0_0_517), .A2(num_leading_zeros[4]), .ZN(n_0_0_417));
   AOI211_X1 i_0_0_512 (.A(n_0_0_421), .B(n_0_0_418), .C1(n_0_0_420), .C2(
      n_0_0_462), .ZN(Sum[23]));
   NOR2_X1 i_0_0_513 (.A1(n_0_0_462), .A2(n_0_0_419), .ZN(n_0_0_418));
   NAND2_X1 i_0_0_514 (.A1(n_0_0_520), .A2(num_leading_zeros[0]), .ZN(n_0_0_419));
   NOR2_X1 i_0_0_515 (.A1(num_leading_zeros[0]), .A2(n_0_0_442), .ZN(n_0_0_420));
   NOR2_X1 i_0_0_516 (.A1(n_0_0_520), .A2(exp_Sum[0]), .ZN(n_0_0_421));
   OAI21_X1 i_0_0_517 (.A(n_0_0_424), .B1(n_0_0_422), .B2(n_0_0_442), .ZN(
      Sum[24]));
   XNOR2_X1 i_0_0_518 (.A(n_0_0_460), .B(n_0_0_423), .ZN(n_0_0_422));
   XNOR2_X1 i_0_0_519 (.A(num_leading_zeros[1]), .B(n_0_0_464), .ZN(n_0_0_423));
   NAND2_X1 i_0_0_520 (.A1(exp_Sum[1]), .A2(n_0_0_442), .ZN(n_0_0_424));
   OAI21_X1 i_0_0_521 (.A(n_0_0_427), .B1(n_0_0_425), .B2(n_0_0_442), .ZN(
      Sum[25]));
   XNOR2_X1 i_0_0_522 (.A(n_0_0_457), .B(n_0_0_426), .ZN(n_0_0_425));
   XNOR2_X1 i_0_0_523 (.A(num_leading_zeros[2]), .B(n_0_0_455), .ZN(n_0_0_426));
   NAND2_X1 i_0_0_524 (.A1(exp_Sum[2]), .A2(n_0_0_442), .ZN(n_0_0_427));
   OAI21_X1 i_0_0_525 (.A(n_0_0_430), .B1(n_0_0_428), .B2(n_0_0_442), .ZN(
      Sum[26]));
   XNOR2_X1 i_0_0_526 (.A(n_0_0_452), .B(n_0_0_429), .ZN(n_0_0_428));
   XNOR2_X1 i_0_0_527 (.A(n_0_0_517), .B(n_0_0_466), .ZN(n_0_0_429));
   NAND2_X1 i_0_0_528 (.A1(exp_Sum[3]), .A2(n_0_0_442), .ZN(n_0_0_430));
   OAI21_X1 i_0_0_529 (.A(n_0_0_433), .B1(n_0_0_431), .B2(n_0_0_442), .ZN(
      Sum[27]));
   XNOR2_X1 i_0_0_530 (.A(n_0_0_449), .B(n_0_0_432), .ZN(n_0_0_431));
   XNOR2_X1 i_0_0_531 (.A(num_leading_zeros[4]), .B(n_0_0_471), .ZN(n_0_0_432));
   NAND2_X1 i_0_0_532 (.A1(exp_Sum[4]), .A2(n_0_0_442), .ZN(n_0_0_433));
   AOI21_X1 i_0_0_533 (.A(n_0_0_434), .B1(n_0_0_435), .B2(n_0_0_520), .ZN(
      Sum[28]));
   NOR2_X1 i_0_0_534 (.A1(n_0_0_520), .A2(exp_Sum[5]), .ZN(n_0_0_434));
   XNOR2_X1 i_0_0_535 (.A(n_0_0_447), .B(n_0_0_445), .ZN(n_0_0_435));
   AOI21_X1 i_0_0_536 (.A(n_0_0_437), .B1(n_0_0_436), .B2(n_0_0_520), .ZN(
      Sum[29]));
   XOR2_X1 i_0_0_537 (.A(n_0_0_443), .B(n_0_0_440), .Z(n_0_0_436));
   NOR2_X1 i_0_0_538 (.A1(n_0_0_520), .A2(exp_Sum[6]), .ZN(n_0_0_437));
   XOR2_X1 i_0_0_539 (.A(n_0_0_473), .B(n_0_0_438), .Z(Sum[30]));
   AOI21_X1 i_0_0_540 (.A(n_0_0_439), .B1(n_0_0_442), .B2(n_0_0_6), .ZN(
      n_0_0_438));
   NOR3_X1 i_0_0_541 (.A1(n_0_0_443), .A2(n_0_0_442), .A3(n_0_0_440), .ZN(
      n_0_0_439));
   OAI21_X1 i_0_0_542 (.A(n_0_0_441), .B1(n_0_96), .B2(n_0_0_503), .ZN(n_0_0_440));
   NAND2_X1 i_0_0_543 (.A1(n_0_96), .A2(B[29]), .ZN(n_0_0_441));
   XNOR2_X1 i_0_0_544 (.A(B[31]), .B(A[31]), .ZN(n_0_0_442));
   NAND2_X1 i_0_0_545 (.A1(n_0_0_447), .A2(n_0_0_444), .ZN(n_0_0_443));
   INV_X1 i_0_0_546 (.A(n_0_0_445), .ZN(n_0_0_444));
   OAI21_X1 i_0_0_547 (.A(n_0_0_446), .B1(n_0_96), .B2(n_0_0_502), .ZN(n_0_0_445));
   NAND2_X1 i_0_0_548 (.A1(n_0_96), .A2(B[28]), .ZN(n_0_0_446));
   OAI21_X1 i_0_0_549 (.A(n_0_0_448), .B1(n_0_0_471), .B2(n_0_0_518), .ZN(
      n_0_0_447));
   OR2_X1 i_0_0_550 (.A1(n_0_0_470), .A2(n_0_0_449), .ZN(n_0_0_448));
   AOI21_X1 i_0_0_551 (.A(n_0_0_450), .B1(n_0_0_467), .B2(num_leading_zeros[3]), 
      .ZN(n_0_0_449));
   INV_X1 i_0_0_552 (.A(n_0_0_451), .ZN(n_0_0_450));
   OAI21_X1 i_0_0_553 (.A(n_0_0_452), .B1(n_0_0_467), .B2(num_leading_zeros[3]), 
      .ZN(n_0_0_451));
   OR2_X1 i_0_0_554 (.A1(n_0_0_454), .A2(n_0_0_453), .ZN(n_0_0_452));
   NOR2_X1 i_0_0_555 (.A1(n_0_0_516), .A2(n_0_0_455), .ZN(n_0_0_453));
   AOI21_X1 i_0_0_556 (.A(n_0_0_457), .B1(n_0_0_455), .B2(n_0_0_516), .ZN(
      n_0_0_454));
   OAI21_X1 i_0_0_557 (.A(n_0_0_456), .B1(n_0_96), .B2(n_0_0_500), .ZN(n_0_0_455));
   NAND2_X1 i_0_0_558 (.A1(n_0_96), .A2(B[25]), .ZN(n_0_0_456));
   AOI21_X1 i_0_0_559 (.A(n_0_0_458), .B1(n_0_0_459), .B2(num_leading_zeros[1]), 
      .ZN(n_0_0_457));
   NOR2_X1 i_0_0_560 (.A1(n_0_0_460), .A2(n_0_0_464), .ZN(n_0_0_458));
   NAND2_X1 i_0_0_561 (.A1(n_0_0_460), .A2(n_0_0_464), .ZN(n_0_0_459));
   NOR2_X1 i_0_0_562 (.A1(num_leading_zeros[0]), .A2(n_0_0_461), .ZN(n_0_0_460));
   INV_X1 i_0_0_563 (.A(n_0_0_462), .ZN(n_0_0_461));
   OAI21_X1 i_0_0_564 (.A(n_0_0_463), .B1(n_0_0_474), .B2(n_0_0_511), .ZN(
      n_0_0_462));
   NAND2_X1 i_0_0_565 (.A1(A[23]), .A2(n_0_0_474), .ZN(n_0_0_463));
   OAI21_X1 i_0_0_566 (.A(n_0_0_465), .B1(n_0_0_474), .B2(n_0_0_512), .ZN(
      n_0_0_464));
   NAND2_X1 i_0_0_567 (.A1(A[24]), .A2(n_0_0_474), .ZN(n_0_0_465));
   INV_X1 i_0_0_568 (.A(n_0_0_467), .ZN(n_0_0_466));
   AND2_X1 i_0_0_569 (.A1(n_0_0_469), .A2(n_0_0_468), .ZN(n_0_0_467));
   NAND2_X1 i_0_0_570 (.A1(n_0_96), .A2(B[26]), .ZN(n_0_0_468));
   NAND2_X1 i_0_0_571 (.A1(A[26]), .A2(n_0_0_474), .ZN(n_0_0_469));
   AND2_X1 i_0_0_572 (.A1(n_0_0_518), .A2(n_0_0_471), .ZN(n_0_0_470));
   OAI21_X1 i_0_0_573 (.A(n_0_0_472), .B1(n_0_96), .B2(n_0_0_501), .ZN(n_0_0_471));
   NAND2_X1 i_0_0_574 (.A1(n_0_96), .A2(B[27]), .ZN(n_0_0_472));
   NOR2_X1 i_0_0_575 (.A1(B[30]), .A2(A[30]), .ZN(n_0_0_473));
   MUX2_X1 i_0_0_576 (.A(A[31]), .B(B[31]), .S(n_0_96), .Z(Sum[31]));
   INV_X1 i_0_0_577 (.A(n_0_0_474), .ZN(n_0_96));
   AOI21_X1 i_0_0_578 (.A(n_0_0_475), .B1(n_0_0_504), .B2(B[30]), .ZN(n_0_0_474));
   NOR2_X1 i_0_0_579 (.A1(n_0_0_477), .A2(n_0_0_476), .ZN(n_0_0_475));
   NOR2_X1 i_0_0_580 (.A1(n_0_0_504), .A2(B[30]), .ZN(n_0_0_476));
   AOI21_X1 i_0_0_581 (.A(n_0_0_483), .B1(n_0_0_478), .B2(n_0_0_480), .ZN(
      n_0_0_477));
   OAI21_X1 i_0_0_582 (.A(n_0_0_482), .B1(n_0_0_484), .B2(n_0_0_479), .ZN(
      n_0_0_478));
   NOR2_X1 i_0_0_583 (.A1(n_0_0_502), .A2(B[28]), .ZN(n_0_0_479));
   NAND2_X1 i_0_0_584 (.A1(n_0_0_514), .A2(A[29]), .ZN(n_0_0_480));
   NOR2_X1 i_0_0_585 (.A1(n_0_0_503), .A2(B[29]), .ZN(n_0_0_481));
   NAND2_X1 i_0_0_586 (.A1(n_0_0_502), .A2(B[28]), .ZN(n_0_0_482));
   NOR2_X1 i_0_0_587 (.A1(n_0_0_514), .A2(A[29]), .ZN(n_0_0_483));
   OAI21_X1 i_0_0_588 (.A(n_0_0_485), .B1(n_0_0_501), .B2(B[27]), .ZN(n_0_0_484));
   NAND2_X1 i_0_0_589 (.A1(n_0_0_487), .A2(n_0_0_486), .ZN(n_0_0_485));
   NAND2_X1 i_0_0_590 (.A1(n_0_0_501), .A2(B[27]), .ZN(n_0_0_486));
   AOI21_X1 i_0_0_591 (.A(n_0_0_488), .B1(n_0_0_491), .B2(n_0_0_489), .ZN(
      n_0_0_487));
   NOR2_X1 i_0_0_592 (.A1(n_0_0_513), .A2(A[26]), .ZN(n_0_0_488));
   NAND2_X1 i_0_0_593 (.A1(n_0_0_513), .A2(A[26]), .ZN(n_0_0_489));
   NOR2_X1 i_0_0_594 (.A1(n_0_0_501), .A2(B[27]), .ZN(n_0_0_490));
   OAI21_X1 i_0_0_595 (.A(n_0_0_492), .B1(n_0_0_493), .B2(n_0_0_495), .ZN(
      n_0_0_491));
   NAND2_X1 i_0_0_596 (.A1(n_0_0_500), .A2(B[25]), .ZN(n_0_0_492));
   AOI21_X1 i_0_0_597 (.A(n_0_0_494), .B1(n_0_0_496), .B2(n_0_0_497), .ZN(
      n_0_0_493));
   NOR2_X1 i_0_0_598 (.A1(n_0_0_512), .A2(A[24]), .ZN(n_0_0_494));
   NOR2_X1 i_0_0_599 (.A1(n_0_0_500), .A2(B[25]), .ZN(n_0_0_495));
   NAND2_X1 i_0_0_600 (.A1(n_0_0_512), .A2(A[24]), .ZN(n_0_0_496));
   NAND2_X1 i_0_0_601 (.A1(n_0_0_511), .A2(A[23]), .ZN(n_0_0_497));
   INV_X1 i_0_0_602 (.A(A[2]), .ZN(n_0_0_498));
   INV_X1 i_0_0_603 (.A(A[21]), .ZN(n_0_0_499));
   INV_X1 i_0_0_604 (.A(A[25]), .ZN(n_0_0_500));
   INV_X1 i_0_0_605 (.A(A[27]), .ZN(n_0_0_501));
   INV_X1 i_0_0_606 (.A(A[28]), .ZN(n_0_0_502));
   INV_X1 i_0_0_607 (.A(A[29]), .ZN(n_0_0_503));
   INV_X1 i_0_0_608 (.A(A[30]), .ZN(n_0_0_504));
   INV_X1 i_0_0_609 (.A(B[17]), .ZN(n_0_0_505));
   INV_X1 i_0_0_610 (.A(B[18]), .ZN(n_0_0_506));
   INV_X1 i_0_0_611 (.A(B[19]), .ZN(n_0_0_507));
   INV_X1 i_0_0_612 (.A(B[20]), .ZN(n_0_0_508));
   INV_X1 i_0_0_613 (.A(B[21]), .ZN(n_0_0_509));
   INV_X1 i_0_0_614 (.A(B[22]), .ZN(n_0_0_510));
   INV_X1 i_0_0_615 (.A(B[23]), .ZN(n_0_0_511));
   INV_X1 i_0_0_616 (.A(B[24]), .ZN(n_0_0_512));
   INV_X1 i_0_0_617 (.A(B[26]), .ZN(n_0_0_513));
   INV_X1 i_0_0_618 (.A(B[29]), .ZN(n_0_0_514));
   INV_X1 i_0_0_619 (.A(n_0_1), .ZN(n_0_0_515));
   INV_X1 i_0_0_620 (.A(num_leading_zeros[2]), .ZN(n_0_0_516));
   INV_X1 i_0_0_621 (.A(num_leading_zeros[3]), .ZN(n_0_0_517));
   INV_X1 i_0_0_622 (.A(num_leading_zeros[4]), .ZN(n_0_0_518));
   INV_X1 i_0_0_623 (.A(n_0_0_482), .ZN(n_0_0_519));
   INV_X1 i_0_0_624 (.A(n_0_0_442), .ZN(n_0_0_520));
   INV_X1 i_0_0_625 (.A(n_0_0_149), .ZN(n_0_0_521));
   INV_X1 i_0_0_626 (.A(n_0_0_310), .ZN(n_0_0_522));
   INV_X1 i_0_0_627 (.A(n_0_0_313), .ZN(n_0_0_523));
   INV_X1 i_0_0_628 (.A(n_0_0_419), .ZN(n_0_0_524));
   INV_X1 i_0_0_629 (.A(n_0_0_420), .ZN(n_0_0_525));
   INV_X1 i_0_0_630 (.A(n_0_0_387), .ZN(n_0_0_526));
   INV_X1 i_0_0_631 (.A(n_0_0_388), .ZN(n_0_0_527));
endmodule
