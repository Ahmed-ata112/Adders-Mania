
// 	Sun Dec  4 17:25:44 2022
//	vlsi
//	localhost.localdomain

module registerNbits (clk, reset, en, inp, out);

output [7:0] out;
input clk;
input en;
input [7:0] inp;
input reset;
wire n_0_0;
wire n_1;
wire n_0;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;


AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk), .E (n_1), .SE (1'b0 ));

endmodule //registerNbits

module registerNbits__0_9 (clk, reset, en, inp, out);

output [7:0] out;
input clk;
input en;
input [7:0] inp;
input reset;
wire n_0_1;
wire n_1;
wire n_0;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;


AND2_X1 i_0_9 (.ZN (n_9), .A1 (inp[7]), .A2 (n_0_1));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (inp[6]), .A2 (n_0_1));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (inp[5]), .A2 (n_0_1));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (inp[4]), .A2 (n_0_1));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (inp[3]), .A2 (n_0_1));
INV_X1 i_0_1 (.ZN (n_0_1), .A (reset));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_1), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_1), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_1), .A2 (inp[0]));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk), .E (n_1), .SE (1'b0 ));

endmodule //registerNbits__0_9

module datapath (inputB, inputA, result);

output [15:0] result;
input [7:0] inputA;
input [7:0] inputB;
wire n_51;
wire n_404;
wire n_405;
wire n_403;
wire n_397;
wire n_43;
wire n_42;
wire n_40;
wire n_2;
wire n_277;
wire n_3;
wire n_338;
wire n_4;
wire n_423;
wire n_424;
wire n_421;
wire n_5;
wire n_339;
wire n_6;
wire n_14;
wire n_7;
wire n_31;
wire n_37;
wire n_30;
wire n_8;
wire n_11;
wire n_36;
wire n_343;
wire n_10;
wire n_9;
wire n_33;
wire n_35;
wire n_12;
wire n_15;
wire n_13;
wire n_255;
wire n_21;
wire n_378;
wire n_60;
wire n_17;
wire n_16;
wire n_18;
wire n_246;
wire n_243;
wire n_244;
wire n_19;
wire n_20;
wire n_22;
wire n_23;
wire n_248;
wire n_24;
wire n_25;
wire n_26;
wire n_230;
wire n_227;
wire n_27;
wire n_228;
wire n_28;
wire n_29;
wire n_32;
wire n_34;
wire n_0;
wire n_157;
wire n_151;
wire n_1;
wire n_65;
wire n_379;
wire n_381;
wire n_380;
wire n_38;
wire n_39;
wire n_41;
wire n_377;
wire n_44;
wire n_45;
wire n_46;
wire n_47;
wire n_48;
wire n_49;
wire n_52;
wire n_50;
wire n_58;
wire n_57;
wire n_54;
wire n_53;
wire n_56;
wire n_59;
wire n_55;
wire n_61;
wire n_62;
wire n_63;
wire n_64;
wire n_67;
wire n_68;
wire n_69;
wire n_70;
wire n_71;
wire n_72;
wire n_73;
wire n_74;
wire n_75;
wire n_76;
wire n_77;
wire n_96;
wire n_78;
wire n_80;
wire n_79;
wire n_83;
wire n_81;
wire n_88;
wire n_82;
wire n_85;
wire n_84;
wire n_89;
wire n_90;
wire n_86;
wire n_87;
wire n_98;
wire n_92;
wire n_91;
wire n_94;
wire n_93;
wire n_95;
wire n_102;
wire n_100;
wire n_104;
wire n_103;
wire n_107;
wire n_110;
wire n_108;
wire n_132;
wire n_105;
wire n_106;
wire n_115;
wire n_109;
wire n_111;
wire n_114;
wire n_112;
wire n_124;
wire n_134;
wire n_125;
wire n_113;
wire n_133;
wire n_122;
wire n_116;
wire n_119;
wire n_117;
wire n_118;
wire n_121;
wire n_120;
wire n_123;
wire n_131;
wire n_126;
wire n_128;
wire n_127;
wire n_129;
wire n_130;
wire n_135;
wire n_136;
wire n_137;
wire n_138;
wire n_139;
wire n_140;
wire n_141;
wire n_142;
wire n_143;
wire n_144;
wire n_145;
wire n_146;
wire n_147;
wire n_148;
wire n_149;
wire n_150;
wire n_154;
wire n_155;
wire n_156;
wire n_159;
wire n_160;
wire n_161;
wire n_162;
wire n_163;
wire n_164;
wire n_165;
wire n_166;
wire n_167;
wire n_168;
wire n_169;
wire n_170;
wire n_171;
wire n_172;
wire n_173;
wire n_174;
wire n_175;
wire n_176;
wire n_177;
wire n_178;
wire n_179;
wire n_180;
wire n_181;
wire n_182;
wire n_183;
wire n_184;
wire n_185;
wire n_186;
wire n_187;
wire n_188;
wire n_189;
wire n_190;
wire n_257;
wire n_258;
wire n_191;
wire n_192;
wire n_193;
wire n_194;
wire n_195;
wire n_196;
wire n_197;
wire n_198;
wire n_199;
wire n_200;
wire n_201;
wire n_202;
wire n_203;
wire n_204;
wire n_205;
wire n_206;
wire n_207;
wire n_209;
wire n_208;
wire n_251;
wire n_211;
wire n_210;
wire n_214;
wire n_212;
wire n_213;
wire n_234;
wire n_250;
wire n_236;
wire n_215;
wire n_218;
wire n_216;
wire n_219;
wire n_217;
wire n_225;
wire n_231;
wire n_226;
wire n_252;
wire n_221;
wire n_220;
wire n_223;
wire n_222;
wire n_224;
wire n_229;
wire n_253;
wire n_385;
wire n_233;
wire n_232;
wire n_412;
wire n_413;
wire n_235;
wire n_249;
wire n_237;
wire n_247;
wire n_238;
wire n_240;
wire n_256;
wire n_242;
wire n_241;
wire n_245;
wire n_254;
wire n_291;
wire n_259;
wire n_261;
wire n_260;
wire n_263;
wire n_262;
wire n_264;
wire n_265;
wire n_275;
wire n_266;
wire n_269;
wire n_267;
wire n_270;
wire n_273;
wire n_271;
wire n_268;
wire n_272;
wire n_274;
wire n_285;
wire n_276;
wire n_278;
wire n_283;
wire n_279;
wire n_281;
wire n_280;
wire n_282;
wire n_284;
wire n_287;
wire n_286;
wire n_290;
wire n_289;
wire n_288;
wire n_410;
wire n_416;
wire n_292;
wire n_293;
wire n_294;
wire n_295;
wire n_297;
wire n_315;
wire n_299;
wire n_301;
wire n_300;
wire n_303;
wire n_302;
wire n_305;
wire n_304;
wire n_313;
wire n_311;
wire n_306;
wire n_307;
wire n_314;
wire n_310;
wire n_309;
wire n_308;
wire n_336;
wire n_337;
wire n_409;
wire n_316;
wire n_312;
wire n_318;
wire n_317;
wire n_320;
wire n_319;
wire n_346;
wire n_340;
wire n_321;
wire n_334;
wire n_322;
wire n_324;
wire n_323;
wire n_330;
wire n_325;
wire n_326;
wire n_332;
wire n_329;
wire n_327;
wire n_328;
wire n_344;
wire n_333;
wire n_342;
wire n_331;
wire n_422;
wire n_426;
wire n_335;
wire n_345;
wire n_341;
wire n_420;
wire n_347;
wire n_348;
wire n_349;
wire n_350;
wire n_351;
wire n_352;
wire n_353;
wire n_354;
wire n_355;
wire n_356;
wire n_357;
wire n_358;
wire n_359;
wire n_360;
wire n_361;
wire n_363;
wire n_364;
wire n_365;
wire n_366;
wire n_367;
wire n_368;
wire n_369;
wire n_370;
wire n_371;
wire n_372;
wire n_373;
wire n_374;
wire n_375;
wire n_376;
wire n_382;
wire n_383;
wire n_384;
wire n_386;
wire n_387;
wire n_388;
wire n_389;
wire n_390;
wire n_391;
wire n_392;
wire n_393;
wire n_394;
wire n_395;
wire n_396;
wire n_398;
wire n_401;
wire n_402;
wire n_399;
wire n_400;
wire n_407;
wire n_406;
wire n_408;
wire n_411;
wire n_414;
wire n_417;
wire n_419;
wire n_418;
wire n_425;


AND2_X1 i_438 (.ZN (n_426), .A1 (inputB[7]), .A2 (inputA[4]));
NAND2_X1 i_437 (.ZN (n_425), .A1 (inputB[5]), .A2 (inputA[5]));
NAND4_X1 i_436 (.ZN (n_424), .A1 (inputB[5]), .A2 (inputA[5]), .A3 (inputB[4]), .A4 (inputA[6]));
NAND2_X1 i_435 (.ZN (n_423), .A1 (inputB[6]), .A2 (inputA[4]));
NAND2_X1 i_434 (.ZN (n_422), .A1 (n_424), .A2 (n_423));
OAI21_X1 i_433 (.ZN (n_421), .A (n_425), .B1 (n_377), .B2 (n_100));
AOI21_X1 i_432 (.ZN (n_420), .A (n_426), .B1 (n_422), .B2 (n_421));
NAND2_X1 i_431 (.ZN (n_419), .A1 (n_413), .A2 (n_233));
NAND2_X1 i_430 (.ZN (n_418), .A1 (n_222), .A2 (n_221));
AOI22_X1 i_427 (.ZN (n_417), .A1 (n_412), .A2 (n_419), .B1 (n_223), .B2 (n_418));
INV_X1 i_426 (.ZN (n_416), .A (n_417));
NAND2_X1 i_423 (.ZN (n_414), .A1 (inputB[4]), .A2 (inputA[4]));
NAND4_X1 i_421 (.ZN (n_413), .A1 (inputB[4]), .A2 (inputA[4]), .A3 (inputB[3]), .A4 (inputA[5]));
OAI21_X1 i_418 (.ZN (n_412), .A (n_414), .B1 (n_159), .B2 (n_65));
AOI22_X1 i_417 (.ZN (n_411), .A1 (n_233), .A2 (n_413), .B1 (n_222), .B2 (n_221));
NAND3_X1 i_416 (.ZN (n_410), .A1 (n_412), .A2 (n_411), .A3 (n_223));
NAND2_X1 i_415 (.ZN (n_409), .A1 (n_288), .A2 (n_410));
INV_X1 i_414 (.ZN (n_408), .A (n_386));
AOI21_X1 i_413 (.ZN (n_407), .A (n_408), .B1 (n_384), .B2 (n_387));
INV_X1 i_412 (.ZN (n_406), .A (n_407));
OAI21_X1 i_411 (.ZN (n_405), .A (n_406), .B1 (n_385), .B2 (n_378));
NAND3_X1 i_410 (.ZN (n_404), .A1 (inputB[7]), .A2 (n_407), .A3 (inputA[7]));
AOI21_X1 i_409 (.ZN (n_403), .A (n_392), .B1 (n_376), .B2 (n_395));
AND2_X1 i_408 (.ZN (n_402), .A1 (n_405), .A2 (n_404));
OAI21_X1 i_407 (.ZN (n_401), .A (n_402), .B1 (n_397), .B2 (n_403));
OAI21_X1 i_406 (.ZN (n_400), .A (n_393), .B1 (n_369), .B2 (n_375));
NAND2_X1 i_405 (.ZN (n_399), .A1 (n_391), .A2 (n_400));
OAI21_X1 i_404 (.ZN (n_398), .A (n_401), .B1 (n_402), .B2 (n_399));
INV_X1 i_403 (.ZN (result[14]), .A (n_398));
INV_X1 i_402 (.ZN (n_397), .A (n_391));
XNOR2_X1 i_401 (.ZN (result[13]), .A (n_394), .B (n_396));
NAND2_X1 i_400 (.ZN (n_396), .A1 (n_376), .A2 (n_395));
INV_X1 i_399 (.ZN (n_395), .A (n_369));
NAND2_X1 i_398 (.ZN (n_394), .A1 (n_393), .A2 (n_391));
INV_X1 i_397 (.ZN (n_393), .A (n_392));
NOR2_X1 i_395 (.ZN (n_392), .A1 (n_389), .A2 (n_390));
NAND2_X1 i_394 (.ZN (n_391), .A1 (n_389), .A2 (n_390));
OAI21_X1 i_393 (.ZN (n_390), .A (n_366), .B1 (n_353), .B2 (n_348));
XOR2_X1 i_392 (.Z (n_389), .A (n_384), .B (n_388));
NAND2_X1 i_391 (.ZN (n_388), .A1 (n_386), .A2 (n_387));
NAND4_X1 i_390 (.ZN (n_387), .A1 (inputA[6]), .A2 (inputB[7]), .A3 (inputA[7]), .A4 (inputB[6]));
OAI22_X1 i_389 (.ZN (n_386), .A1 (n_377), .A2 (n_385), .B1 (n_378), .B2 (n_255));
INV_X1 i_388 (.ZN (n_385), .A (inputB[7]));
OAI21_X1 i_387 (.ZN (n_384), .A (n_379), .B1 (n_382), .B2 (n_383));
INV_X1 i_386 (.ZN (n_383), .A (n_381));
INV_X1 i_385 (.ZN (n_382), .A (n_380));
NAND2_X1 i_384 (.ZN (n_381), .A1 (inputA[5]), .A2 (inputB[7]));
NAND4_X1 i_383 (.ZN (n_380), .A1 (inputB[5]), .A2 (inputA[6]), .A3 (inputA[7]), .A4 (inputB[6]));
OAI22_X1 i_382 (.ZN (n_379), .A1 (n_377), .A2 (n_255), .B1 (n_378), .B2 (n_157));
INV_X1 i_381 (.ZN (n_378), .A (inputA[7]));
INV_X1 i_380 (.ZN (n_377), .A (inputA[6]));
INV_X1 i_379 (.ZN (n_376), .A (n_375));
AOI21_X1 i_378 (.ZN (n_375), .A (n_370), .B1 (n_373), .B2 (n_374));
NAND3_X1 i_377 (.ZN (n_374), .A1 (n_300), .A2 (n_261), .A3 (n_319));
AOI221_X1 i_376 (.ZN (n_373), .A (n_371), .B1 (n_340), .B2 (n_321), .C1 (n_372), .C2 (n_305));
AND3_X1 i_374 (.ZN (n_372), .A1 (n_319), .A2 (n_303), .A3 (n_304));
INV_X1 i_373 (.ZN (n_371), .A (n_360));
INV_X1 i_372 (.ZN (n_370), .A (n_359));
NOR3_X1 i_370 (.ZN (n_369), .A1 (n_367), .A2 (n_368), .A3 (n_260));
INV_X1 i_369 (.ZN (n_368), .A (n_211));
NAND4_X1 i_368 (.ZN (n_367), .A1 (n_292), .A2 (n_300), .A3 (n_319), .A4 (n_359));
INV_X1 i_367 (.ZN (n_366), .A (n_354));
XNOR2_X1 i_366 (.ZN (result[12]), .A (n_361), .B (n_365));
OAI21_X1 i_365 (.ZN (n_365), .A (n_320), .B1 (n_363), .B2 (n_364));
NAND2_X1 i_364 (.ZN (n_364), .A1 (n_300), .A2 (n_319));
NOR2_X1 i_363 (.ZN (n_363), .A1 (n_299), .A2 (n_315));
NAND2_X1 i_361 (.ZN (n_361), .A1 (n_359), .A2 (n_360));
NAND2_X1 i_360 (.ZN (n_360), .A1 (n_356), .A2 (n_358));
OR2_X1 i_359 (.ZN (n_359), .A1 (n_356), .A2 (n_358));
AND2_X1 i_358 (.ZN (n_358), .A1 (n_357), .A2 (n_324));
NAND2_X1 i_357 (.ZN (n_357), .A1 (n_323), .A2 (n_334));
XNOR2_X1 i_356 (.ZN (n_356), .A (n_355), .B (n_348));
NOR2_X1 i_355 (.ZN (n_355), .A1 (n_353), .A2 (n_354));
NOR2_X1 i_354 (.ZN (n_354), .A1 (n_351), .A2 (n_352));
AND2_X1 i_353 (.ZN (n_353), .A1 (n_351), .A2 (n_352));
OAI21_X1 i_352 (.ZN (n_352), .A (n_43), .B1 (n_41), .B2 (n_39));
NOR2_X1 i_351 (.ZN (n_351), .A1 (n_349), .A2 (n_350));
INV_X1 i_350 (.ZN (n_350), .A (n_38));
AOI21_X1 i_349 (.ZN (n_349), .A (n_381), .B1 (n_379), .B2 (n_380));
OAI21_X1 i_348 (.ZN (n_348), .A (n_344), .B1 (n_347), .B2 (n_332));
INV_X1 i_347 (.ZN (n_347), .A (n_333));
INV_X1 i_346 (.ZN (n_346), .A (n_301));
INV_X1 i_345 (.ZN (n_345), .A (n_5));
INV_X1 i_344 (.ZN (n_344), .A (n_420));
INV_X1 i_343 (.ZN (n_343), .A (n_37));
INV_X1 i_342 (.ZN (n_342), .A (n_2));
NAND2_X1 i_341 (.ZN (n_341), .A1 (n_313), .A2 (n_306));
NAND2_X1 i_340 (.ZN (n_340), .A1 (n_311), .A2 (n_341));
OAI21_X1 i_339 (.ZN (n_339), .A (n_15), .B1 (n_7), .B2 (n_16));
NAND3_X1 i_338 (.ZN (n_338), .A1 (n_421), .A2 (n_424), .A3 (n_423));
NAND3_X1 i_337 (.ZN (n_337), .A1 (n_345), .A2 (n_338), .A3 (n_339));
OAI21_X1 i_335 (.ZN (n_336), .A (n_6), .B1 (n_5), .B2 (n_4));
INV_X1 i_334 (.ZN (n_335), .A (n_336));
OAI21_X1 i_333 (.ZN (n_334), .A (n_337), .B1 (n_309), .B2 (n_335));
NAND3_X1 i_332 (.ZN (n_333), .A1 (n_422), .A2 (n_426), .A3 (n_421));
AOI21_X1 i_331 (.ZN (n_332), .A (n_343), .B1 (n_31), .B2 (n_30));
AOI21_X1 i_330 (.ZN (n_331), .A (n_42), .B1 (n_43), .B2 (n_40));
NOR2_X1 i_329 (.ZN (n_330), .A1 (n_342), .A2 (n_331));
NAND2_X1 i_328 (.ZN (n_329), .A1 (n_344), .A2 (n_333));
AOI21_X1 i_327 (.ZN (n_328), .A (n_10), .B1 (n_11), .B2 (n_36));
INV_X1 i_326 (.ZN (n_327), .A (n_328));
AOI21_X1 i_325 (.ZN (n_326), .A (n_329), .B1 (n_37), .B2 (n_327));
AOI21_X1 i_324 (.ZN (n_325), .A (n_326), .B1 (n_332), .B2 (n_329));
NAND2_X1 i_323 (.ZN (n_324), .A1 (n_330), .A2 (n_325));
OR2_X1 i_322 (.ZN (n_323), .A1 (n_330), .A2 (n_325));
NAND2_X1 i_321 (.ZN (n_322), .A1 (n_324), .A2 (n_323));
XOR2_X1 i_320 (.Z (n_321), .A (n_334), .B (n_322));
NAND2_X1 i_319 (.ZN (n_320), .A1 (n_340), .A2 (n_321));
OR2_X1 i_318 (.ZN (n_319), .A1 (n_340), .A2 (n_321));
OAI21_X1 i_317 (.ZN (n_318), .A (n_300), .B1 (n_346), .B2 (n_315));
NAND2_X1 i_316 (.ZN (n_317), .A1 (n_320), .A2 (n_319));
XOR2_X1 i_315 (.Z (result[11]), .A (n_318), .B (n_317));
INV_X1 i_314 (.ZN (n_316), .A (n_278));
AOI21_X1 i_313 (.ZN (n_315), .A (n_260), .B1 (n_291), .B2 (n_262));
AOI221_X1 i_312 (.ZN (n_314), .A (n_316), .B1 (n_285), .B2 (n_277), .C1 (n_409), .C2 (n_416));
INV_X1 i_311 (.ZN (n_313), .A (n_314));
AOI21_X1 i_310 (.ZN (n_312), .A (n_3), .B1 (n_287), .B2 (n_286));
OAI211_X1 i_309 (.ZN (n_311), .A (n_409), .B (n_416), .C1 (n_316), .C2 (n_312));
INV_X1 i_308 (.ZN (n_310), .A (n_311));
NAND2_X1 i_307 (.ZN (n_309), .A1 (n_8), .A2 (n_9));
NAND2_X1 i_306 (.ZN (n_308), .A1 (n_336), .A2 (n_337));
XOR2_X1 i_305 (.Z (n_307), .A (n_309), .B (n_308));
INV_X1 i_304 (.ZN (n_306), .A (n_307));
OAI21_X1 i_303 (.ZN (n_305), .A (n_307), .B1 (n_314), .B2 (n_310));
NAND3_X1 i_302 (.ZN (n_304), .A1 (n_313), .A2 (n_311), .A3 (n_306));
OAI21_X1 i_301 (.ZN (n_303), .A (n_267), .B1 (n_270), .B2 (n_275));
AND2_X1 i_300 (.ZN (n_302), .A1 (n_305), .A2 (n_304));
NAND2_X1 i_299 (.ZN (n_301), .A1 (n_303), .A2 (n_302));
OR2_X1 i_298 (.ZN (n_300), .A1 (n_303), .A2 (n_302));
NAND2_X1 i_297 (.ZN (n_299), .A1 (n_301), .A2 (n_300));
XNOR2_X1 i_295 (.ZN (result[10]), .A (n_315), .B (n_299));
INV_X1 i_294 (.ZN (n_297), .A (n_173));
NAND3_X1 i_292 (.ZN (n_295), .A1 (n_173), .A2 (n_105), .A3 (n_104));
OAI211_X1 i_291 (.ZN (n_294), .A (n_174), .B (n_295), .C1 (n_106), .C2 (n_297));
NAND2_X1 i_290 (.ZN (n_293), .A1 (n_206), .A2 (n_294));
NAND3_X1 i_289 (.ZN (n_292), .A1 (n_210), .A2 (n_293), .A3 (n_205));
NAND2_X1 i_288 (.ZN (n_291), .A1 (n_211), .A2 (n_292));
NAND2_X1 i_287 (.ZN (n_290), .A1 (n_410), .A2 (n_416));
AOI21_X1 i_286 (.ZN (n_289), .A (n_240), .B1 (n_241), .B2 (n_247));
INV_X1 i_285 (.ZN (n_288), .A (n_289));
NAND2_X1 i_284 (.ZN (n_287), .A1 (n_290), .A2 (n_289));
OR2_X1 i_283 (.ZN (n_286), .A1 (n_290), .A2 (n_289));
NAND2_X1 i_282 (.ZN (n_285), .A1 (n_287), .A2 (n_286));
AND3_X1 i_281 (.ZN (n_284), .A1 (n_17), .A2 (n_14), .A3 (n_15));
AOI21_X1 i_280 (.ZN (n_283), .A (n_284), .B1 (n_13), .B2 (n_16));
OAI21_X1 i_279 (.ZN (n_282), .A (n_34), .B1 (n_12), .B2 (n_32));
INV_X1 i_278 (.ZN (n_281), .A (n_282));
AND3_X1 i_277 (.ZN (n_280), .A1 (n_35), .A2 (n_33), .A3 (n_36));
NOR2_X1 i_276 (.ZN (n_279), .A1 (n_281), .A2 (n_280));
OR2_X1 i_275 (.ZN (n_278), .A1 (n_283), .A2 (n_279));
NAND2_X1 i_274 (.ZN (n_277), .A1 (n_283), .A2 (n_279));
NAND2_X1 i_273 (.ZN (n_276), .A1 (n_278), .A2 (n_277));
XOR2_X1 i_272 (.Z (n_275), .A (n_285), .B (n_276));
NOR2_X1 i_271 (.ZN (n_274), .A1 (n_231), .A2 (n_226));
OAI21_X1 i_270 (.ZN (n_273), .A (n_225), .B1 (n_219), .B2 (n_274));
OAI21_X1 i_269 (.ZN (n_272), .A (n_254), .B1 (n_250), .B2 (n_236));
NAND2_X1 i_268 (.ZN (n_271), .A1 (n_234), .A2 (n_272));
NOR2_X1 i_267 (.ZN (n_270), .A1 (n_273), .A2 (n_271));
INV_X1 i_266 (.ZN (n_269), .A (n_270));
AOI21_X1 i_265 (.ZN (n_268), .A (n_196), .B1 (n_249), .B2 (n_237));
OAI21_X1 i_264 (.ZN (n_267), .A (n_273), .B1 (n_235), .B2 (n_268));
AOI21_X1 i_263 (.ZN (n_266), .A (n_270), .B1 (n_273), .B2 (n_271));
AOI21_X1 i_262 (.ZN (n_265), .A (n_275), .B1 (n_269), .B2 (n_267));
AOI21_X1 i_261 (.ZN (n_264), .A (n_265), .B1 (n_275), .B2 (n_266));
INV_X1 i_260 (.ZN (n_263), .A (n_264));
NAND2_X1 i_259 (.ZN (n_262), .A1 (n_215), .A2 (n_263));
INV_X1 i_258 (.ZN (n_261), .A (n_262));
NOR2_X1 i_257 (.ZN (n_260), .A1 (n_215), .A2 (n_263));
NOR2_X1 i_256 (.ZN (n_259), .A1 (n_261), .A2 (n_260));
XNOR2_X1 i_255 (.ZN (result[9]), .A (n_291), .B (n_259));
INV_X1 i_254 (.ZN (n_258), .A (n_23));
INV_X1 i_253 (.ZN (n_257), .A (n_26));
INV_X1 i_252 (.ZN (n_256), .A (n_18));
INV_X1 i_251 (.ZN (n_255), .A (inputB[6]));
INV_X1 i_250 (.ZN (n_254), .A (n_196));
INV_X1 i_249 (.ZN (n_253), .A (n_155));
INV_X1 i_248 (.ZN (n_252), .A (n_198));
INV_X1 i_247 (.ZN (n_251), .A (n_206));
OAI21_X1 i_246 (.ZN (n_250), .A (n_187), .B1 (n_186), .B2 (n_180));
INV_X1 i_245 (.ZN (n_249), .A (n_250));
OAI21_X1 i_244 (.ZN (n_248), .A (n_25), .B1 (n_157), .B2 (n_67));
OAI21_X1 i_243 (.ZN (n_247), .A (n_248), .B1 (n_258), .B2 (n_257));
OAI21_X1 i_242 (.ZN (n_246), .A (n_20), .B1 (n_100), .B2 (n_21));
INV_X1 i_241 (.ZN (n_245), .A (n_246));
NAND4_X1 i_240 (.ZN (n_244), .A1 (inputB[4]), .A2 (inputB[3]), .A3 (inputA[4]), .A4 (inputA[3]));
NAND2_X1 i_239 (.ZN (n_243), .A1 (inputB[2]), .A2 (inputA[5]));
AOI21_X1 i_238 (.ZN (n_242), .A (n_245), .B1 (n_244), .B2 (n_243));
NAND2_X1 i_237 (.ZN (n_241), .A1 (n_256), .A2 (n_242));
NOR2_X1 i_236 (.ZN (n_240), .A1 (n_256), .A2 (n_242));
AOI21_X1 i_234 (.ZN (n_238), .A (n_240), .B1 (n_256), .B2 (n_242));
XOR2_X1 i_233 (.Z (n_237), .A (n_247), .B (n_238));
INV_X1 i_232 (.ZN (n_236), .A (n_237));
NOR2_X1 i_231 (.ZN (n_235), .A1 (n_249), .A2 (n_237));
INV_X1 i_230 (.ZN (n_234), .A (n_235));
NAND2_X1 i_229 (.ZN (n_233), .A1 (inputB[5]), .A2 (inputA[3]));
NAND2_X1 i_228 (.ZN (n_232), .A1 (n_412), .A2 (n_413));
XOR2_X1 i_227 (.Z (n_231), .A (n_233), .B (n_232));
OAI21_X1 i_226 (.ZN (n_230), .A (n_29), .B1 (n_385), .B2 (n_45));
INV_X1 i_225 (.ZN (n_229), .A (n_230));
OAI21_X1 i_224 (.ZN (n_228), .A (n_154), .B1 (n_253), .B2 (n_150));
NAND4_X1 i_223 (.ZN (n_227), .A1 (inputB[7]), .A2 (inputB[0]), .A3 (inputA[7]), .A4 (inputA[0]));
AOI21_X1 i_222 (.ZN (n_226), .A (n_229), .B1 (n_228), .B2 (n_227));
NAND2_X1 i_221 (.ZN (n_225), .A1 (n_231), .A2 (n_226));
NAND2_X1 i_220 (.ZN (n_224), .A1 (inputB[2]), .A2 (inputA[6]));
OAI21_X1 i_219 (.ZN (n_223), .A (n_224), .B1 (n_67), .B2 (n_255));
NAND4_X1 i_218 (.ZN (n_222), .A1 (inputB[2]), .A2 (inputA[6]), .A3 (inputB[6]), .A4 (inputA[2]));
NAND2_X1 i_217 (.ZN (n_221), .A1 (inputB[1]), .A2 (inputA[7]));
NAND2_X1 i_216 (.ZN (n_220), .A1 (n_223), .A2 (n_222));
XNOR2_X1 i_215 (.ZN (n_219), .A (n_221), .B (n_220));
AOI21_X1 i_214 (.ZN (n_218), .A (n_252), .B1 (n_199), .B2 (n_202));
OAI21_X1 i_213 (.ZN (n_217), .A (n_225), .B1 (n_231), .B2 (n_226));
XNOR2_X1 i_212 (.ZN (n_216), .A (n_219), .B (n_217));
NOR2_X1 i_211 (.ZN (n_215), .A1 (n_218), .A2 (n_216));
AOI21_X1 i_210 (.ZN (n_214), .A (n_215), .B1 (n_218), .B2 (n_216));
OAI21_X1 i_209 (.ZN (n_213), .A (n_234), .B1 (n_250), .B2 (n_236));
XOR2_X1 i_208 (.Z (n_212), .A (n_196), .B (n_213));
OR2_X1 i_207 (.ZN (n_211), .A1 (n_214), .A2 (n_212));
NAND2_X1 i_206 (.ZN (n_210), .A1 (n_214), .A2 (n_212));
NAND2_X1 i_205 (.ZN (n_209), .A1 (n_211), .A2 (n_210));
AOI21_X1 i_204 (.ZN (n_208), .A (n_251), .B1 (n_205), .B2 (n_177));
XNOR2_X1 i_203 (.ZN (result[8]), .A (n_209), .B (n_208));
XOR2_X1 i_202 (.Z (result[7]), .A (n_207), .B (n_177));
NAND2_X1 i_201 (.ZN (n_207), .A1 (n_205), .A2 (n_206));
NAND2_X1 i_200 (.ZN (n_206), .A1 (n_203), .A2 (n_142));
NAND3_X1 i_199 (.ZN (n_205), .A1 (n_204), .A2 (n_137), .A3 (n_139));
INV_X1 i_198 (.ZN (n_204), .A (n_203));
XOR2_X1 i_197 (.Z (n_203), .A (n_200), .B (n_202));
NAND2_X1 i_196 (.ZN (n_202), .A1 (n_201), .A2 (n_167));
NAND2_X1 i_195 (.ZN (n_201), .A1 (n_170), .A2 (n_166));
NAND2_X1 i_194 (.ZN (n_200), .A1 (n_198), .A2 (n_199));
NAND2_X1 i_193 (.ZN (n_199), .A1 (n_189), .A2 (n_197));
OR2_X1 i_192 (.ZN (n_198), .A1 (n_189), .A2 (n_197));
OAI21_X1 i_191 (.ZN (n_197), .A (n_196), .B1 (n_192), .B2 (n_195));
NAND2_X1 i_190 (.ZN (n_196), .A1 (n_192), .A2 (n_195));
NAND2_X1 i_189 (.ZN (n_195), .A1 (n_193), .A2 (n_194));
NAND2_X1 i_188 (.ZN (n_194), .A1 (n_28), .A2 (n_27));
NAND3_X1 i_187 (.ZN (n_193), .A1 (n_230), .A2 (n_227), .A3 (n_228));
NAND2_X1 i_186 (.ZN (n_192), .A1 (n_190), .A2 (n_191));
OAI21_X1 i_185 (.ZN (n_191), .A (n_257), .B1 (n_24), .B2 (n_258));
NAND3_X1 i_184 (.ZN (n_190), .A1 (n_26), .A2 (n_23), .A3 (n_248));
XNOR2_X1 i_183 (.ZN (n_189), .A (n_188), .B (n_180));
NAND2_X1 i_182 (.ZN (n_188), .A1 (n_187), .A2 (n_185));
OR2_X1 i_181 (.ZN (n_187), .A1 (n_182), .A2 (n_184));
INV_X1 i_180 (.ZN (n_186), .A (n_185));
NAND2_X1 i_179 (.ZN (n_185), .A1 (n_182), .A2 (n_184));
OAI21_X1 i_178 (.ZN (n_184), .A (n_160), .B1 (n_183), .B2 (n_156));
INV_X1 i_177 (.ZN (n_183), .A (n_161));
NAND2_X1 i_176 (.ZN (n_182), .A1 (n_181), .A2 (n_149));
NAND2_X1 i_175 (.ZN (n_181), .A1 (n_146), .A2 (n_143));
NOR2_X1 i_174 (.ZN (n_180), .A1 (n_178), .A2 (n_179));
INV_X1 i_173 (.ZN (n_179), .A (n_19));
AOI21_X1 i_172 (.ZN (n_178), .A (n_243), .B1 (n_246), .B2 (n_244));
OAI21_X1 i_171 (.ZN (n_177), .A (n_173), .B1 (n_176), .B2 (n_136));
INV_X1 i_170 (.ZN (n_176), .A (n_174));
XNOR2_X1 i_169 (.ZN (result[6]), .A (n_175), .B (n_136));
NAND2_X1 i_168 (.ZN (n_175), .A1 (n_173), .A2 (n_174));
NAND2_X1 i_167 (.ZN (n_174), .A1 (n_171), .A2 (n_172));
OR2_X1 i_166 (.ZN (n_173), .A1 (n_171), .A2 (n_172));
AOI21_X1 i_165 (.ZN (n_172), .A (n_141), .B1 (n_124), .B2 (n_140));
XNOR2_X1 i_164 (.ZN (n_171), .A (n_168), .B (n_170));
XOR2_X1 i_163 (.Z (n_170), .A (n_169), .B (n_143));
NAND2_X1 i_162 (.ZN (n_169), .A1 (n_146), .A2 (n_149));
NAND2_X1 i_161 (.ZN (n_168), .A1 (n_166), .A2 (n_167));
NAND2_X1 i_160 (.ZN (n_167), .A1 (n_163), .A2 (n_165));
OR2_X1 i_159 (.ZN (n_166), .A1 (n_163), .A2 (n_165));
XNOR2_X1 i_158 (.ZN (n_165), .A (n_164), .B (n_156));
NAND2_X1 i_157 (.ZN (n_164), .A1 (n_160), .A2 (n_161));
XNOR2_X1 i_156 (.ZN (n_163), .A (n_162), .B (n_150));
NAND2_X1 i_155 (.ZN (n_162), .A1 (n_154), .A2 (n_155));
NAND4_X1 i_154 (.ZN (n_161), .A1 (inputB[1]), .A2 (inputA[5]), .A3 (inputB[5]), .A4 (inputA[1]));
OAI22_X1 i_153 (.ZN (n_160), .A1 (n_44), .A2 (n_159), .B1 (n_157), .B2 (n_59));
INV_X1 i_152 (.ZN (n_159), .A (inputA[5]));
INV_X1 i_150 (.ZN (n_157), .A (inputB[5]));
AND2_X1 i_149 (.ZN (n_156), .A1 (inputB[0]), .A2 (inputA[6]));
NAND4_X1 i_148 (.ZN (n_155), .A1 (inputB[3]), .A2 (inputA[3]), .A3 (inputB[2]), .A4 (inputA[4]));
OAI22_X1 i_147 (.ZN (n_154), .A1 (n_65), .A2 (n_21), .B1 (n_151), .B2 (n_60));
INV_X1 i_142 (.ZN (n_151), .A (inputA[4]));
AND2_X1 i_141 (.ZN (n_150), .A1 (inputB[4]), .A2 (inputA[2]));
OAI21_X1 i_139 (.ZN (n_149), .A (n_144), .B1 (n_147), .B2 (n_148));
INV_X1 i_138 (.ZN (n_148), .A (n_119));
AND2_X1 i_137 (.ZN (n_147), .A1 (n_117), .A2 (n_123));
OAI211_X1 i_136 (.ZN (n_146), .A (n_145), .B (n_119), .C1 (n_118), .C2 (n_122));
INV_X1 i_135 (.ZN (n_145), .A (n_144));
NAND2_X1 i_134 (.ZN (n_144), .A1 (inputB[6]), .A2 (inputA[0]));
OAI21_X1 i_132 (.ZN (n_143), .A (n_129), .B1 (n_127), .B2 (n_130));
INV_X1 i_131 (.ZN (n_142), .A (n_141));
NOR2_X1 i_130 (.ZN (n_141), .A1 (n_140), .A2 (n_124));
INV_X1 i_129 (.ZN (n_140), .A (n_139));
NAND2_X1 i_128 (.ZN (n_139), .A1 (n_138), .A2 (n_111));
OAI21_X1 i_127 (.ZN (n_138), .A (n_115), .B1 (n_114), .B2 (n_112));
INV_X1 i_126 (.ZN (n_137), .A (n_124));
NAND2_X1 i_125 (.ZN (n_136), .A1 (n_135), .A2 (n_106));
NAND2_X1 i_124 (.ZN (n_135), .A1 (n_104), .A2 (n_105));
INV_X1 i_123 (.ZN (n_134), .A (n_89));
INV_X1 i_122 (.ZN (n_133), .A (n_93));
INV_X1 i_121 (.ZN (n_132), .A (n_80));
NAND2_X1 i_120 (.ZN (n_131), .A1 (inputB[5]), .A2 (inputA[0]));
INV_X1 i_119 (.ZN (n_130), .A (n_131));
OAI21_X1 i_118 (.ZN (n_129), .A (n_22), .B1 (n_100), .B2 (n_59));
INV_X1 i_117 (.ZN (n_128), .A (n_129));
AND4_X1 i_116 (.ZN (n_127), .A1 (inputB[4]), .A2 (inputB[0]), .A3 (inputA[5]), .A4 (inputA[1]));
NOR2_X1 i_115 (.ZN (n_126), .A1 (n_128), .A2 (n_127));
XNOR2_X1 i_114 (.ZN (n_125), .A (n_131), .B (n_126));
NAND3_X1 i_113 (.ZN (n_124), .A1 (n_90), .A2 (n_125), .A3 (n_72));
NAND2_X1 i_112 (.ZN (n_123), .A1 (inputB[1]), .A2 (inputA[4]));
INV_X1 i_111 (.ZN (n_122), .A (n_123));
NAND2_X1 i_110 (.ZN (n_121), .A1 (inputB[2]), .A2 (inputA[3]));
NAND2_X1 i_109 (.ZN (n_120), .A1 (inputB[3]), .A2 (inputA[2]));
NAND2_X1 i_108 (.ZN (n_119), .A1 (n_121), .A2 (n_120));
NOR2_X1 i_107 (.ZN (n_118), .A1 (n_121), .A2 (n_120));
INV_X1 i_106 (.ZN (n_117), .A (n_118));
NAND2_X1 i_105 (.ZN (n_116), .A1 (n_119), .A2 (n_117));
XNOR2_X1 i_104 (.ZN (n_115), .A (n_122), .B (n_116));
AOI21_X1 i_103 (.ZN (n_114), .A (n_86), .B1 (n_87), .B2 (n_84));
OAI21_X1 i_102 (.ZN (n_113), .A (n_94), .B1 (n_133), .B2 (n_92));
INV_X1 i_101 (.ZN (n_112), .A (n_113));
NAND2_X1 i_100 (.ZN (n_111), .A1 (n_114), .A2 (n_112));
OAI21_X1 i_99 (.ZN (n_110), .A (n_124), .B1 (n_134), .B2 (n_125));
OAI21_X1 i_98 (.ZN (n_109), .A (n_111), .B1 (n_114), .B2 (n_112));
XOR2_X1 i_97 (.Z (n_108), .A (n_115), .B (n_109));
NOR2_X1 i_96 (.ZN (n_107), .A1 (n_110), .A2 (n_108));
INV_X1 i_95 (.ZN (n_106), .A (n_107));
NAND2_X1 i_94 (.ZN (n_105), .A1 (n_110), .A2 (n_108));
AOI21_X1 i_93 (.ZN (n_104), .A (n_132), .B1 (n_79), .B2 (n_95));
AOI21_X1 i_92 (.ZN (n_103), .A (n_107), .B1 (n_110), .B2 (n_108));
XOR2_X1 i_91 (.Z (result[5]), .A (n_104), .B (n_103));
INV_X1 i_90 (.ZN (n_102), .A (n_75));
INV_X1 i_88 (.ZN (n_100), .A (inputB[4]));
INV_X1 i_86 (.ZN (n_98), .A (n_68));
AOI21_X1 i_84 (.ZN (n_96), .A (n_102), .B1 (n_76), .B2 (n_62));
INV_X1 i_83 (.ZN (n_95), .A (n_96));
OAI22_X1 i_82 (.ZN (n_94), .A1 (n_65), .A2 (n_59), .B1 (n_67), .B2 (n_60));
NAND4_X1 i_81 (.ZN (n_93), .A1 (inputB[3]), .A2 (inputB[2]), .A3 (inputA[2]), .A4 (inputA[1]));
AND2_X1 i_80 (.ZN (n_92), .A1 (inputA[3]), .A2 (inputB[1]));
NAND2_X1 i_79 (.ZN (n_91), .A1 (n_94), .A2 (n_93));
XNOR2_X1 i_78 (.ZN (n_90), .A (n_92), .B (n_91));
NAND2_X1 i_77 (.ZN (n_89), .A1 (n_72), .A2 (n_90));
AOI21_X1 i_76 (.ZN (n_88), .A (n_98), .B1 (n_69), .B2 (n_64));
INV_X1 i_75 (.ZN (n_87), .A (n_88));
AOI22_X1 i_74 (.ZN (n_86), .A1 (inputA[4]), .A2 (inputB[0]), .B1 (inputB[4]), .B2 (inputA[0]));
INV_X1 i_73 (.ZN (n_85), .A (n_86));
NAND4_X1 i_72 (.ZN (n_84), .A1 (inputA[4]), .A2 (inputB[0]), .A3 (inputA[0]), .A4 (inputB[4]));
OAI21_X1 i_71 (.ZN (n_83), .A (n_89), .B1 (n_72), .B2 (n_90));
NAND2_X1 i_70 (.ZN (n_82), .A1 (n_85), .A2 (n_84));
XOR2_X1 i_69 (.Z (n_81), .A (n_88), .B (n_82));
NAND2_X1 i_68 (.ZN (n_80), .A1 (n_83), .A2 (n_81));
OR2_X1 i_67 (.ZN (n_79), .A1 (n_83), .A2 (n_81));
NAND2_X1 i_66 (.ZN (n_78), .A1 (n_80), .A2 (n_79));
XNOR2_X1 i_65 (.ZN (result[4]), .A (n_96), .B (n_78));
XOR2_X1 i_64 (.Z (result[3]), .A (n_77), .B (n_62));
NAND2_X1 i_63 (.ZN (n_77), .A1 (n_75), .A2 (n_76));
NAND2_X1 i_62 (.ZN (n_76), .A1 (n_71), .A2 (n_74));
OR2_X1 i_61 (.ZN (n_75), .A1 (n_71), .A2 (n_74));
AOI21_X1 i_60 (.ZN (n_74), .A (n_72), .B1 (n_54), .B2 (n_73));
NAND2_X1 i_59 (.ZN (n_73), .A1 (inputB[0]), .A2 (inputA[3]));
INV_X1 i_58 (.ZN (n_72), .A (n_63));
XOR2_X1 i_57 (.Z (n_71), .A (n_70), .B (n_64));
NAND2_X1 i_56 (.ZN (n_70), .A1 (n_68), .A2 (n_69));
NAND4_X1 i_55 (.ZN (n_69), .A1 (inputB[1]), .A2 (inputA[2]), .A3 (inputB[3]), .A4 (inputA[0]));
OAI22_X1 i_54 (.ZN (n_68), .A1 (n_44), .A2 (n_67), .B1 (n_65), .B2 (n_45));
INV_X1 i_53 (.ZN (n_67), .A (inputA[2]));
INV_X1 i_51 (.ZN (n_65), .A (inputB[3]));
NAND2_X1 i_50 (.ZN (n_64), .A1 (inputB[2]), .A2 (inputA[1]));
NAND4_X1 i_49 (.ZN (n_63), .A1 (n_55), .A2 (inputA[3]), .A3 (inputA[1]), .A4 (inputB[1]));
OAI21_X1 i_48 (.ZN (n_62), .A (n_57), .B1 (n_61), .B2 (n_52));
INV_X1 i_47 (.ZN (n_61), .A (n_58));
INV_X1 i_46 (.ZN (n_60), .A (inputB[2]));
INV_X1 i_45 (.ZN (n_59), .A (inputA[1]));
OR2_X1 i_44 (.ZN (n_58), .A1 (n_49), .A2 (n_60));
OAI21_X1 i_43 (.ZN (n_57), .A (n_49), .B1 (n_60), .B2 (n_45));
NAND2_X1 i_42 (.ZN (n_56), .A1 (inputB[0]), .A2 (inputA[2]));
INV_X1 i_41 (.ZN (n_55), .A (n_56));
NAND3_X1 i_40 (.ZN (n_54), .A1 (inputB[1]), .A2 (n_55), .A3 (inputA[1]));
OAI21_X1 i_39 (.ZN (n_53), .A (n_56), .B1 (n_59), .B2 (n_44));
AND2_X1 i_38 (.ZN (n_52), .A1 (n_54), .A2 (n_53));
NAND2_X1 i_37 (.ZN (n_50), .A1 (n_58), .A2 (n_57));
XNOR2_X1 i_36 (.ZN (result[2]), .A (n_52), .B (n_50));
AOI21_X1 i_35 (.ZN (result[1]), .A (n_48), .B1 (n_46), .B2 (n_47));
INV_X1 i_34 (.ZN (n_49), .A (n_48));
NOR2_X1 i_33 (.ZN (n_48), .A1 (n_46), .A2 (n_47));
NAND2_X1 i_32 (.ZN (n_47), .A1 (inputB[1]), .A2 (inputA[0]));
NAND2_X1 i_31 (.ZN (n_46), .A1 (inputB[0]), .A2 (inputA[1]));
INV_X1 i_30 (.ZN (n_45), .A (inputA[0]));
INV_X1 i_29 (.ZN (n_44), .A (inputB[1]));
AND2_X1 i_28 (.ZN (result[0]), .A1 (inputB[0]), .A2 (inputA[0]));
OAI22_X1 i_27 (.ZN (n_43), .A1 (n_157), .A2 (n_377), .B1 (n_255), .B2 (n_159));
NAND2_X1 i_26 (.ZN (n_42), .A1 (inputA[7]), .A2 (inputB[4]));
INV_X1 i_508 (.ZN (n_41), .A (n_42));
NAND4_X1 i_25 (.ZN (n_40), .A1 (inputB[6]), .A2 (inputB[5]), .A3 (inputA[6]), .A4 (inputA[5]));
INV_X1 i_506 (.ZN (n_39), .A (n_40));
NAND3_X1 i_502 (.ZN (n_38), .A1 (n_379), .A2 (n_381), .A3 (n_380));
NAND2_X1 i_24 (.ZN (n_1), .A1 (inputB[7]), .A2 (inputA[3]));
OAI21_X1 i_23 (.ZN (n_37), .A (n_1), .B1 (n_378), .B2 (n_65));
NAND2_X1 i_22 (.ZN (n_0), .A1 (inputB[4]), .A2 (inputA[5]));
OAI21_X1 i_21 (.ZN (n_36), .A (n_0), .B1 (n_157), .B2 (n_151));
NAND2_X1 i_20 (.ZN (n_35), .A1 (inputA[6]), .A2 (inputB[3]));
INV_X1 i_19 (.ZN (n_34), .A (n_35));
NAND4_X1 i_18 (.ZN (n_33), .A1 (inputB[5]), .A2 (inputB[4]), .A3 (inputA[5]), .A4 (inputA[4]));
INV_X1 i_17 (.ZN (n_32), .A (n_33));
OAI21_X1 i_16 (.ZN (n_31), .A (n_36), .B1 (n_32), .B2 (n_34));
NAND4_X1 i_15 (.ZN (n_30), .A1 (inputB[7]), .A2 (inputB[3]), .A3 (inputA[7]), .A4 (inputA[3]));
NAND2_X1 i_463 (.ZN (n_29), .A1 (inputA[7]), .A2 (inputB[0]));
INV_X1 i_429 (.ZN (n_28), .A (n_228));
NAND2_X1 i_428 (.ZN (n_27), .A1 (n_230), .A2 (n_227));
NAND2_X1 i_424 (.ZN (n_26), .A1 (inputB[6]), .A2 (inputA[1]));
NAND2_X1 i_422 (.ZN (n_25), .A1 (inputA[6]), .A2 (inputB[1]));
INV_X1 i_420 (.ZN (n_24), .A (n_248));
NAND4_X1 i_419 (.ZN (n_23), .A1 (inputB[5]), .A2 (inputB[1]), .A3 (inputA[6]), .A4 (inputA[2]));
NAND2_X1 i_396 (.ZN (n_22), .A1 (inputA[5]), .A2 (inputB[0]));
INV_X1 i_14 (.ZN (n_21), .A (inputA[3]));
NAND2_X1 i_375 (.ZN (n_20), .A1 (inputB[3]), .A2 (inputA[4]));
NAND3_X1 i_371 (.ZN (n_19), .A1 (n_246), .A2 (n_243), .A3 (n_244));
NAND2_X1 i_336 (.ZN (n_18), .A1 (inputB[7]), .A2 (inputA[1]));
NAND2_X1 i_13 (.ZN (n_17), .A1 (inputB[7]), .A2 (inputA[2]));
INV_X1 i_12 (.ZN (n_16), .A (n_17));
OAI22_X1 i_11 (.ZN (n_15), .A1 (n_255), .A2 (n_21), .B1 (n_378), .B2 (n_60));
NAND4_X1 i_10 (.ZN (n_14), .A1 (inputB[6]), .A2 (inputB[2]), .A3 (inputA[7]), .A4 (inputA[3]));
NAND2_X1 i_9 (.ZN (n_13), .A1 (n_15), .A2 (n_14));
INV_X1 i_8 (.ZN (n_12), .A (n_36));
NAND2_X1 i_7 (.ZN (n_11), .A1 (n_33), .A2 (n_35));
INV_X1 i_6 (.ZN (n_10), .A (n_30));
OAI211_X1 i_5 (.ZN (n_9), .A (n_11), .B (n_36), .C1 (n_343), .C2 (n_10));
NAND3_X1 i_4 (.ZN (n_8), .A1 (n_31), .A2 (n_37), .A3 (n_30));
INV_X1 i_145 (.ZN (n_7), .A (n_14));
INV_X1 i_143 (.ZN (n_6), .A (n_339));
AOI21_X1 i_3 (.ZN (n_5), .A (n_423), .B1 (n_424), .B2 (n_421));
INV_X1 i_140 (.ZN (n_4), .A (n_338));
INV_X1 i_133 (.ZN (n_3), .A (n_277));
NAND3_X1 i_2 (.ZN (n_2), .A1 (n_43), .A2 (n_42), .A3 (n_40));
OAI21_X1 i_1 (.ZN (n_51), .A (n_405), .B1 (n_403), .B2 (n_397));
NAND2_X1 i_0 (.ZN (result[15]), .A1 (n_51), .A2 (n_404));

endmodule //datapath

module multiplyTimes (inputA, inputB, result);

output [15:0] result;
input [7:0] inputA;
input [7:0] inputB;


datapath i_0 (.result ({result[15], result[14], result[13], result[12], result[11], 
    result[10], result[9], result[8], result[7], result[6], result[5], result[4], 
    result[3], result[2], result[1], result[0]}), .inputA ({inputA[7], inputA[6], 
    inputA[5], inputA[4], inputA[3], inputA[2], inputA[1], inputA[0]}), .inputB ({
    inputB[7], inputB[6], inputB[5], inputB[4], inputB[3], inputB[2], inputB[1], 
    inputB[0]}));

endmodule //multiplyTimes

module registerNbits__0_6 (clk, reset, en, inp, out);

output [7:0] out;
input clk;
input en;
input [7:0] inp;
input reset;
wire n_0_0;
wire n_1;
wire n_0;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;


AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk), .E (n_1), .SE (1'b0 ));

endmodule //registerNbits__0_6

module registerNbits__0_3 (clk, reset, en, inp, out);

output [7:0] out;
input clk;
input en;
input [7:0] inp;
input reset;
wire n_0_0;
wire n_1;
wire n_0;
wire n_9;
wire n_8;
wire n_7;
wire n_6;
wire n_5;
wire n_4;
wire n_3;
wire n_2;


AND2_X1 i_0_9 (.ZN (n_9), .A1 (n_0_0), .A2 (inp[7]));
AND2_X1 i_0_8 (.ZN (n_8), .A1 (n_0_0), .A2 (inp[6]));
AND2_X1 i_0_7 (.ZN (n_7), .A1 (n_0_0), .A2 (inp[5]));
AND2_X1 i_0_6 (.ZN (n_6), .A1 (n_0_0), .A2 (inp[4]));
AND2_X1 i_0_5 (.ZN (n_5), .A1 (n_0_0), .A2 (inp[3]));
AND2_X1 i_0_4 (.ZN (n_4), .A1 (n_0_0), .A2 (inp[2]));
AND2_X1 i_0_3 (.ZN (n_3), .A1 (n_0_0), .A2 (inp[1]));
AND2_X1 i_0_2 (.ZN (n_2), .A1 (n_0_0), .A2 (inp[0]));
INV_X1 i_0_1 (.ZN (n_0_0), .A (reset));
OR2_X1 i_0_0 (.ZN (n_1), .A1 (en), .A2 (reset));
DFF_X1 \out_reg[0]  (.Q (out[0]), .CK (n_0), .D (n_2));
DFF_X1 \out_reg[1]  (.Q (out[1]), .CK (n_0), .D (n_3));
DFF_X1 \out_reg[2]  (.Q (out[2]), .CK (n_0), .D (n_4));
DFF_X1 \out_reg[3]  (.Q (out[3]), .CK (n_0), .D (n_5));
DFF_X1 \out_reg[4]  (.Q (out[4]), .CK (n_0), .D (n_6));
DFF_X1 \out_reg[5]  (.Q (out[5]), .CK (n_0), .D (n_7));
DFF_X1 \out_reg[6]  (.Q (out[6]), .CK (n_0), .D (n_8));
DFF_X1 \out_reg[7]  (.Q (out[7]), .CK (n_0), .D (n_9));
CLKGATETST_X1 clk_gate_out_reg (.GCK (n_0), .CK (clk), .E (n_1), .SE (1'b0 ));

endmodule //registerNbits__0_3

module integrationMult (clk, reset, en, inputA, inputB, result);

output [15:0] result;
input clk;
input en;
input [7:0] inputA;
input [7:0] inputB;
input reset;
wire \A_reg[7] ;
wire \A_reg[6] ;
wire \A_reg[5] ;
wire \A_reg[4] ;
wire \A_reg[3] ;
wire \A_reg[2] ;
wire \A_reg[1] ;
wire \A_reg[0] ;
wire \B_reg[7] ;
wire \B_reg[6] ;
wire \B_reg[5] ;
wire \B_reg[4] ;
wire \B_reg[3] ;
wire \B_reg[2] ;
wire \B_reg[1] ;
wire \B_reg[0] ;
wire \outB_reg[7] ;
wire \outB_reg[6] ;
wire \outB_reg[5] ;
wire \outB_reg[4] ;
wire \outB_reg[3] ;
wire \outB_reg[2] ;
wire \outB_reg[1] ;
wire \outB_reg[0] ;
wire \outA_reg[7] ;
wire \outA_reg[6] ;
wire \outA_reg[5] ;
wire \outA_reg[4] ;
wire \outA_reg[3] ;
wire \outA_reg[2] ;
wire \outA_reg[1] ;
wire \outA_reg[0] ;


registerNbits outA (.out ({result[7], result[6], result[5], result[4], result[3], 
    result[2], result[1], result[0]}), .clk (clk), .en (en), .inp ({\outB_reg[7] , 
    \outB_reg[6] , \outB_reg[5] , \outB_reg[4] , \outB_reg[3] , \outB_reg[2] , \outB_reg[1] , 
    \outB_reg[0] }), .reset (reset));
registerNbits__0_9 outB (.out ({result[15], result[14], result[13], result[12], result[11], 
    result[10], result[9], result[8]}), .clk (clk), .en (en), .inp ({\outA_reg[7] , 
    \outA_reg[6] , \outA_reg[5] , \outA_reg[4] , \outA_reg[3] , \outA_reg[2] , \outA_reg[1] , 
    \outA_reg[0] }), .reset (reset));
multiplyTimes mult (.result ({\outA_reg[7] , \outA_reg[6] , \outA_reg[5] , \outA_reg[4] , 
    \outA_reg[3] , \outA_reg[2] , \outA_reg[1] , \outA_reg[0] , \outB_reg[7] , \outB_reg[6] , 
    \outB_reg[5] , \outB_reg[4] , \outB_reg[3] , \outB_reg[2] , \outB_reg[1] , \outB_reg[0] })
    , .inputA ({\A_reg[7] , \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , \A_reg[2] , 
    \A_reg[1] , \A_reg[0] }), .inputB ({\B_reg[7] , \B_reg[6] , \B_reg[5] , \B_reg[4] , 
    \B_reg[3] , \B_reg[2] , \B_reg[1] , \B_reg[0] }));
registerNbits__0_6 regB (.out ({\B_reg[7] , \B_reg[6] , \B_reg[5] , \B_reg[4] , \B_reg[3] , 
    \B_reg[2] , \B_reg[1] , \B_reg[0] }), .clk (clk), .en (en), .inp ({inputB[7], 
    inputB[6], inputB[5], inputB[4], inputB[3], inputB[2], inputB[1], inputB[0]}), .reset (reset));
registerNbits__0_3 regA (.out ({\A_reg[7] , \A_reg[6] , \A_reg[5] , \A_reg[4] , \A_reg[3] , 
    \A_reg[2] , \A_reg[1] , \A_reg[0] }), .clk (clk), .en (en), .inp ({inputA[7], 
    inputA[6], inputA[5], inputA[4], inputA[3], inputA[2], inputA[1], inputA[0]}), .reset (reset));

endmodule //integrationMult


