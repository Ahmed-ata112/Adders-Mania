/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Thu Oct 27 15:15:12 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1109461611 */

module full_adder__0_69(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(o_sum));
   AND2_X1 i_0_1 (.A1(i_bit2), .A2(i_bit1), .ZN(o_carry));
endmodule

module full_adder__0_73(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_77(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_81(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_85(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_89(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_93(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_97(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_101(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_105(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_109(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_113(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_117(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_121(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_125(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_129(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_133(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_137(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_141(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_145(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_149(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_153(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_157(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_161(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_165(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_169(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_173(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_177(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_181(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_185(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_189(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_193(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_197(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_201(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_205(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_209(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_213(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_217(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_221(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_225(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_229(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_233(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_237(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_241(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_245(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_249(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_253(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_257(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_261(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_265(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_269(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_273(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_277(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_281(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_285(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_289(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_293(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_297(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_301(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_305(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_309(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_313(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder__0_317(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module full_adder(i_bit1, i_bit2, i_carry, o_sum, o_carry);
   input i_bit1;
   input i_bit2;
   input i_carry;
   output o_sum;
   output o_carry;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(i_bit1), .B(i_bit2), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(i_carry), .Z(o_sum));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(i_carry), .B1(i_bit1), .B2(i_bit2), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(o_carry));
endmodule

module ripple_adder(i_add1, i_add2, o_result);
   input [63:0]i_add1;
   input [63:0]i_add2;
   output [64:0]o_result;

   full_adder__0_69 genblk1_0_full_adder_inst (.i_bit1(i_add1[0]), .i_bit2(
      i_add2[0]), .i_carry(), .o_sum(o_result[0]), .o_carry(n_0));
   full_adder__0_73 genblk1_1_full_adder_inst (.i_bit1(i_add1[1]), .i_bit2(
      i_add2[1]), .i_carry(n_0), .o_sum(o_result[1]), .o_carry(n_1));
   full_adder__0_77 genblk1_2_full_adder_inst (.i_bit1(i_add1[2]), .i_bit2(
      i_add2[2]), .i_carry(n_1), .o_sum(o_result[2]), .o_carry(n_2));
   full_adder__0_81 genblk1_3_full_adder_inst (.i_bit1(i_add1[3]), .i_bit2(
      i_add2[3]), .i_carry(n_2), .o_sum(o_result[3]), .o_carry(n_3));
   full_adder__0_85 genblk1_4_full_adder_inst (.i_bit1(i_add1[4]), .i_bit2(
      i_add2[4]), .i_carry(n_3), .o_sum(o_result[4]), .o_carry(n_4));
   full_adder__0_89 genblk1_5_full_adder_inst (.i_bit1(i_add1[5]), .i_bit2(
      i_add2[5]), .i_carry(n_4), .o_sum(o_result[5]), .o_carry(n_5));
   full_adder__0_93 genblk1_6_full_adder_inst (.i_bit1(i_add1[6]), .i_bit2(
      i_add2[6]), .i_carry(n_5), .o_sum(o_result[6]), .o_carry(n_6));
   full_adder__0_97 genblk1_7_full_adder_inst (.i_bit1(i_add1[7]), .i_bit2(
      i_add2[7]), .i_carry(n_6), .o_sum(o_result[7]), .o_carry(n_7));
   full_adder__0_101 genblk1_8_full_adder_inst (.i_bit1(i_add1[8]), .i_bit2(
      i_add2[8]), .i_carry(n_7), .o_sum(o_result[8]), .o_carry(n_8));
   full_adder__0_105 genblk1_9_full_adder_inst (.i_bit1(i_add1[9]), .i_bit2(
      i_add2[9]), .i_carry(n_8), .o_sum(o_result[9]), .o_carry(n_9));
   full_adder__0_109 genblk1_10_full_adder_inst (.i_bit1(i_add1[10]), .i_bit2(
      i_add2[10]), .i_carry(n_9), .o_sum(o_result[10]), .o_carry(n_10));
   full_adder__0_113 genblk1_11_full_adder_inst (.i_bit1(i_add1[11]), .i_bit2(
      i_add2[11]), .i_carry(n_10), .o_sum(o_result[11]), .o_carry(n_11));
   full_adder__0_117 genblk1_12_full_adder_inst (.i_bit1(i_add1[12]), .i_bit2(
      i_add2[12]), .i_carry(n_11), .o_sum(o_result[12]), .o_carry(n_12));
   full_adder__0_121 genblk1_13_full_adder_inst (.i_bit1(i_add1[13]), .i_bit2(
      i_add2[13]), .i_carry(n_12), .o_sum(o_result[13]), .o_carry(n_13));
   full_adder__0_125 genblk1_14_full_adder_inst (.i_bit1(i_add1[14]), .i_bit2(
      i_add2[14]), .i_carry(n_13), .o_sum(o_result[14]), .o_carry(n_14));
   full_adder__0_129 genblk1_15_full_adder_inst (.i_bit1(i_add1[15]), .i_bit2(
      i_add2[15]), .i_carry(n_14), .o_sum(o_result[15]), .o_carry(n_15));
   full_adder__0_133 genblk1_16_full_adder_inst (.i_bit1(i_add1[16]), .i_bit2(
      i_add2[16]), .i_carry(n_15), .o_sum(o_result[16]), .o_carry(n_16));
   full_adder__0_137 genblk1_17_full_adder_inst (.i_bit1(i_add1[17]), .i_bit2(
      i_add2[17]), .i_carry(n_16), .o_sum(o_result[17]), .o_carry(n_17));
   full_adder__0_141 genblk1_18_full_adder_inst (.i_bit1(i_add1[18]), .i_bit2(
      i_add2[18]), .i_carry(n_17), .o_sum(o_result[18]), .o_carry(n_18));
   full_adder__0_145 genblk1_19_full_adder_inst (.i_bit1(i_add1[19]), .i_bit2(
      i_add2[19]), .i_carry(n_18), .o_sum(o_result[19]), .o_carry(n_19));
   full_adder__0_149 genblk1_20_full_adder_inst (.i_bit1(i_add1[20]), .i_bit2(
      i_add2[20]), .i_carry(n_19), .o_sum(o_result[20]), .o_carry(n_20));
   full_adder__0_153 genblk1_21_full_adder_inst (.i_bit1(i_add1[21]), .i_bit2(
      i_add2[21]), .i_carry(n_20), .o_sum(o_result[21]), .o_carry(n_21));
   full_adder__0_157 genblk1_22_full_adder_inst (.i_bit1(i_add1[22]), .i_bit2(
      i_add2[22]), .i_carry(n_21), .o_sum(o_result[22]), .o_carry(n_22));
   full_adder__0_161 genblk1_23_full_adder_inst (.i_bit1(i_add1[23]), .i_bit2(
      i_add2[23]), .i_carry(n_22), .o_sum(o_result[23]), .o_carry(n_23));
   full_adder__0_165 genblk1_24_full_adder_inst (.i_bit1(i_add1[24]), .i_bit2(
      i_add2[24]), .i_carry(n_23), .o_sum(o_result[24]), .o_carry(n_24));
   full_adder__0_169 genblk1_25_full_adder_inst (.i_bit1(i_add1[25]), .i_bit2(
      i_add2[25]), .i_carry(n_24), .o_sum(o_result[25]), .o_carry(n_25));
   full_adder__0_173 genblk1_26_full_adder_inst (.i_bit1(i_add1[26]), .i_bit2(
      i_add2[26]), .i_carry(n_25), .o_sum(o_result[26]), .o_carry(n_26));
   full_adder__0_177 genblk1_27_full_adder_inst (.i_bit1(i_add1[27]), .i_bit2(
      i_add2[27]), .i_carry(n_26), .o_sum(o_result[27]), .o_carry(n_27));
   full_adder__0_181 genblk1_28_full_adder_inst (.i_bit1(i_add1[28]), .i_bit2(
      i_add2[28]), .i_carry(n_27), .o_sum(o_result[28]), .o_carry(n_28));
   full_adder__0_185 genblk1_29_full_adder_inst (.i_bit1(i_add1[29]), .i_bit2(
      i_add2[29]), .i_carry(n_28), .o_sum(o_result[29]), .o_carry(n_29));
   full_adder__0_189 genblk1_30_full_adder_inst (.i_bit1(i_add1[30]), .i_bit2(
      i_add2[30]), .i_carry(n_29), .o_sum(o_result[30]), .o_carry(n_30));
   full_adder__0_193 genblk1_31_full_adder_inst (.i_bit1(i_add1[31]), .i_bit2(
      i_add2[31]), .i_carry(n_30), .o_sum(o_result[31]), .o_carry(n_31));
   full_adder__0_197 genblk1_32_full_adder_inst (.i_bit1(i_add1[32]), .i_bit2(
      i_add2[32]), .i_carry(n_31), .o_sum(o_result[32]), .o_carry(n_32));
   full_adder__0_201 genblk1_33_full_adder_inst (.i_bit1(i_add1[33]), .i_bit2(
      i_add2[33]), .i_carry(n_32), .o_sum(o_result[33]), .o_carry(n_33));
   full_adder__0_205 genblk1_34_full_adder_inst (.i_bit1(i_add1[34]), .i_bit2(
      i_add2[34]), .i_carry(n_33), .o_sum(o_result[34]), .o_carry(n_34));
   full_adder__0_209 genblk1_35_full_adder_inst (.i_bit1(i_add1[35]), .i_bit2(
      i_add2[35]), .i_carry(n_34), .o_sum(o_result[35]), .o_carry(n_35));
   full_adder__0_213 genblk1_36_full_adder_inst (.i_bit1(i_add1[36]), .i_bit2(
      i_add2[36]), .i_carry(n_35), .o_sum(o_result[36]), .o_carry(n_36));
   full_adder__0_217 genblk1_37_full_adder_inst (.i_bit1(i_add1[37]), .i_bit2(
      i_add2[37]), .i_carry(n_36), .o_sum(o_result[37]), .o_carry(n_37));
   full_adder__0_221 genblk1_38_full_adder_inst (.i_bit1(i_add1[38]), .i_bit2(
      i_add2[38]), .i_carry(n_37), .o_sum(o_result[38]), .o_carry(n_38));
   full_adder__0_225 genblk1_39_full_adder_inst (.i_bit1(i_add1[39]), .i_bit2(
      i_add2[39]), .i_carry(n_38), .o_sum(o_result[39]), .o_carry(n_39));
   full_adder__0_229 genblk1_40_full_adder_inst (.i_bit1(i_add1[40]), .i_bit2(
      i_add2[40]), .i_carry(n_39), .o_sum(o_result[40]), .o_carry(n_40));
   full_adder__0_233 genblk1_41_full_adder_inst (.i_bit1(i_add1[41]), .i_bit2(
      i_add2[41]), .i_carry(n_40), .o_sum(o_result[41]), .o_carry(n_41));
   full_adder__0_237 genblk1_42_full_adder_inst (.i_bit1(i_add1[42]), .i_bit2(
      i_add2[42]), .i_carry(n_41), .o_sum(o_result[42]), .o_carry(n_42));
   full_adder__0_241 genblk1_43_full_adder_inst (.i_bit1(i_add1[43]), .i_bit2(
      i_add2[43]), .i_carry(n_42), .o_sum(o_result[43]), .o_carry(n_43));
   full_adder__0_245 genblk1_44_full_adder_inst (.i_bit1(i_add1[44]), .i_bit2(
      i_add2[44]), .i_carry(n_43), .o_sum(o_result[44]), .o_carry(n_44));
   full_adder__0_249 genblk1_45_full_adder_inst (.i_bit1(i_add1[45]), .i_bit2(
      i_add2[45]), .i_carry(n_44), .o_sum(o_result[45]), .o_carry(n_45));
   full_adder__0_253 genblk1_46_full_adder_inst (.i_bit1(i_add1[46]), .i_bit2(
      i_add2[46]), .i_carry(n_45), .o_sum(o_result[46]), .o_carry(n_46));
   full_adder__0_257 genblk1_47_full_adder_inst (.i_bit1(i_add1[47]), .i_bit2(
      i_add2[47]), .i_carry(n_46), .o_sum(o_result[47]), .o_carry(n_47));
   full_adder__0_261 genblk1_48_full_adder_inst (.i_bit1(i_add1[48]), .i_bit2(
      i_add2[48]), .i_carry(n_47), .o_sum(o_result[48]), .o_carry(n_48));
   full_adder__0_265 genblk1_49_full_adder_inst (.i_bit1(i_add1[49]), .i_bit2(
      i_add2[49]), .i_carry(n_48), .o_sum(o_result[49]), .o_carry(n_49));
   full_adder__0_269 genblk1_50_full_adder_inst (.i_bit1(i_add1[50]), .i_bit2(
      i_add2[50]), .i_carry(n_49), .o_sum(o_result[50]), .o_carry(n_50));
   full_adder__0_273 genblk1_51_full_adder_inst (.i_bit1(i_add1[51]), .i_bit2(
      i_add2[51]), .i_carry(n_50), .o_sum(o_result[51]), .o_carry(n_51));
   full_adder__0_277 genblk1_52_full_adder_inst (.i_bit1(i_add1[52]), .i_bit2(
      i_add2[52]), .i_carry(n_51), .o_sum(o_result[52]), .o_carry(n_52));
   full_adder__0_281 genblk1_53_full_adder_inst (.i_bit1(i_add1[53]), .i_bit2(
      i_add2[53]), .i_carry(n_52), .o_sum(o_result[53]), .o_carry(n_53));
   full_adder__0_285 genblk1_54_full_adder_inst (.i_bit1(i_add1[54]), .i_bit2(
      i_add2[54]), .i_carry(n_53), .o_sum(o_result[54]), .o_carry(n_54));
   full_adder__0_289 genblk1_55_full_adder_inst (.i_bit1(i_add1[55]), .i_bit2(
      i_add2[55]), .i_carry(n_54), .o_sum(o_result[55]), .o_carry(n_55));
   full_adder__0_293 genblk1_56_full_adder_inst (.i_bit1(i_add1[56]), .i_bit2(
      i_add2[56]), .i_carry(n_55), .o_sum(o_result[56]), .o_carry(n_56));
   full_adder__0_297 genblk1_57_full_adder_inst (.i_bit1(i_add1[57]), .i_bit2(
      i_add2[57]), .i_carry(n_56), .o_sum(o_result[57]), .o_carry(n_57));
   full_adder__0_301 genblk1_58_full_adder_inst (.i_bit1(i_add1[58]), .i_bit2(
      i_add2[58]), .i_carry(n_57), .o_sum(o_result[58]), .o_carry(n_58));
   full_adder__0_305 genblk1_59_full_adder_inst (.i_bit1(i_add1[59]), .i_bit2(
      i_add2[59]), .i_carry(n_58), .o_sum(o_result[59]), .o_carry(n_59));
   full_adder__0_309 genblk1_60_full_adder_inst (.i_bit1(i_add1[60]), .i_bit2(
      i_add2[60]), .i_carry(n_59), .o_sum(o_result[60]), .o_carry(n_60));
   full_adder__0_313 genblk1_61_full_adder_inst (.i_bit1(i_add1[61]), .i_bit2(
      i_add2[61]), .i_carry(n_60), .o_sum(o_result[61]), .o_carry(n_61));
   full_adder__0_317 genblk1_62_full_adder_inst (.i_bit1(i_add1[62]), .i_bit2(
      i_add2[62]), .i_carry(n_61), .o_sum(o_result[62]), .o_carry(n_62));
   full_adder genblk1_63_full_adder_inst (.i_bit1(i_add1[63]), .i_bit2(
      i_add2[63]), .i_carry(n_62), .o_sum(o_result[63]), .o_carry(o_result[64]));
endmodule

module Register(write_data, write_enable, clk, rst, MyData);
   input [64:0]write_data;
   input write_enable;
   input clk;
   input rst;
   output [64:0]MyData;

   CLKGATETST_X1 clk_gate_MyData_reg (.CK(clk), .E(write_enable), .SE(1'b0), 
      .GCK(n_0));
   DFFR_X1 \MyData_reg[64]  (.D(write_data[64]), .RN(n_1), .CK(n_0), .Q(
      MyData[64]), .QN());
   INV_X1 i_0_0 (.A(rst), .ZN(n_1));
   DFFR_X1 \MyData_reg[63]  (.D(write_data[63]), .RN(n_1), .CK(n_0), .Q(
      MyData[63]), .QN());
   DFFR_X1 \MyData_reg[62]  (.D(write_data[62]), .RN(n_1), .CK(n_0), .Q(
      MyData[62]), .QN());
   DFFR_X1 \MyData_reg[61]  (.D(write_data[61]), .RN(n_1), .CK(n_0), .Q(
      MyData[61]), .QN());
   DFFR_X1 \MyData_reg[60]  (.D(write_data[60]), .RN(n_1), .CK(n_0), .Q(
      MyData[60]), .QN());
   DFFR_X1 \MyData_reg[59]  (.D(write_data[59]), .RN(n_1), .CK(n_0), .Q(
      MyData[59]), .QN());
   DFFR_X1 \MyData_reg[58]  (.D(write_data[58]), .RN(n_1), .CK(n_0), .Q(
      MyData[58]), .QN());
   DFFR_X1 \MyData_reg[57]  (.D(write_data[57]), .RN(n_1), .CK(n_0), .Q(
      MyData[57]), .QN());
   DFFR_X1 \MyData_reg[56]  (.D(write_data[56]), .RN(n_1), .CK(n_0), .Q(
      MyData[56]), .QN());
   DFFR_X1 \MyData_reg[55]  (.D(write_data[55]), .RN(n_1), .CK(n_0), .Q(
      MyData[55]), .QN());
   DFFR_X1 \MyData_reg[54]  (.D(write_data[54]), .RN(n_1), .CK(n_0), .Q(
      MyData[54]), .QN());
   DFFR_X1 \MyData_reg[53]  (.D(write_data[53]), .RN(n_1), .CK(n_0), .Q(
      MyData[53]), .QN());
   DFFR_X1 \MyData_reg[52]  (.D(write_data[52]), .RN(n_1), .CK(n_0), .Q(
      MyData[52]), .QN());
   DFFR_X1 \MyData_reg[51]  (.D(write_data[51]), .RN(n_1), .CK(n_0), .Q(
      MyData[51]), .QN());
   DFFR_X1 \MyData_reg[50]  (.D(write_data[50]), .RN(n_1), .CK(n_0), .Q(
      MyData[50]), .QN());
   DFFR_X1 \MyData_reg[49]  (.D(write_data[49]), .RN(n_1), .CK(n_0), .Q(
      MyData[49]), .QN());
   DFFR_X1 \MyData_reg[48]  (.D(write_data[48]), .RN(n_1), .CK(n_0), .Q(
      MyData[48]), .QN());
   DFFR_X1 \MyData_reg[47]  (.D(write_data[47]), .RN(n_1), .CK(n_0), .Q(
      MyData[47]), .QN());
   DFFR_X1 \MyData_reg[46]  (.D(write_data[46]), .RN(n_1), .CK(n_0), .Q(
      MyData[46]), .QN());
   DFFR_X1 \MyData_reg[45]  (.D(write_data[45]), .RN(n_1), .CK(n_0), .Q(
      MyData[45]), .QN());
   DFFR_X1 \MyData_reg[44]  (.D(write_data[44]), .RN(n_1), .CK(n_0), .Q(
      MyData[44]), .QN());
   DFFR_X1 \MyData_reg[43]  (.D(write_data[43]), .RN(n_1), .CK(n_0), .Q(
      MyData[43]), .QN());
   DFFR_X1 \MyData_reg[42]  (.D(write_data[42]), .RN(n_1), .CK(n_0), .Q(
      MyData[42]), .QN());
   DFFR_X1 \MyData_reg[41]  (.D(write_data[41]), .RN(n_1), .CK(n_0), .Q(
      MyData[41]), .QN());
   DFFR_X1 \MyData_reg[40]  (.D(write_data[40]), .RN(n_1), .CK(n_0), .Q(
      MyData[40]), .QN());
   DFFR_X1 \MyData_reg[39]  (.D(write_data[39]), .RN(n_1), .CK(n_0), .Q(
      MyData[39]), .QN());
   DFFR_X1 \MyData_reg[38]  (.D(write_data[38]), .RN(n_1), .CK(n_0), .Q(
      MyData[38]), .QN());
   DFFR_X1 \MyData_reg[37]  (.D(write_data[37]), .RN(n_1), .CK(n_0), .Q(
      MyData[37]), .QN());
   DFFR_X1 \MyData_reg[36]  (.D(write_data[36]), .RN(n_1), .CK(n_0), .Q(
      MyData[36]), .QN());
   DFFR_X1 \MyData_reg[35]  (.D(write_data[35]), .RN(n_1), .CK(n_0), .Q(
      MyData[35]), .QN());
   DFFR_X1 \MyData_reg[34]  (.D(write_data[34]), .RN(n_1), .CK(n_0), .Q(
      MyData[34]), .QN());
   DFFR_X1 \MyData_reg[33]  (.D(write_data[33]), .RN(n_1), .CK(n_0), .Q(
      MyData[33]), .QN());
   DFFR_X1 \MyData_reg[32]  (.D(write_data[32]), .RN(n_1), .CK(n_0), .Q(
      MyData[32]), .QN());
   DFFR_X1 \MyData_reg[31]  (.D(write_data[31]), .RN(n_1), .CK(n_0), .Q(
      MyData[31]), .QN());
   DFFR_X1 \MyData_reg[30]  (.D(write_data[30]), .RN(n_1), .CK(n_0), .Q(
      MyData[30]), .QN());
   DFFR_X1 \MyData_reg[29]  (.D(write_data[29]), .RN(n_1), .CK(n_0), .Q(
      MyData[29]), .QN());
   DFFR_X1 \MyData_reg[28]  (.D(write_data[28]), .RN(n_1), .CK(n_0), .Q(
      MyData[28]), .QN());
   DFFR_X1 \MyData_reg[27]  (.D(write_data[27]), .RN(n_1), .CK(n_0), .Q(
      MyData[27]), .QN());
   DFFR_X1 \MyData_reg[26]  (.D(write_data[26]), .RN(n_1), .CK(n_0), .Q(
      MyData[26]), .QN());
   DFFR_X1 \MyData_reg[25]  (.D(write_data[25]), .RN(n_1), .CK(n_0), .Q(
      MyData[25]), .QN());
   DFFR_X1 \MyData_reg[24]  (.D(write_data[24]), .RN(n_1), .CK(n_0), .Q(
      MyData[24]), .QN());
   DFFR_X1 \MyData_reg[23]  (.D(write_data[23]), .RN(n_1), .CK(n_0), .Q(
      MyData[23]), .QN());
   DFFR_X1 \MyData_reg[22]  (.D(write_data[22]), .RN(n_1), .CK(n_0), .Q(
      MyData[22]), .QN());
   DFFR_X1 \MyData_reg[21]  (.D(write_data[21]), .RN(n_1), .CK(n_0), .Q(
      MyData[21]), .QN());
   DFFR_X1 \MyData_reg[20]  (.D(write_data[20]), .RN(n_1), .CK(n_0), .Q(
      MyData[20]), .QN());
   DFFR_X1 \MyData_reg[19]  (.D(write_data[19]), .RN(n_1), .CK(n_0), .Q(
      MyData[19]), .QN());
   DFFR_X1 \MyData_reg[18]  (.D(write_data[18]), .RN(n_1), .CK(n_0), .Q(
      MyData[18]), .QN());
   DFFR_X1 \MyData_reg[17]  (.D(write_data[17]), .RN(n_1), .CK(n_0), .Q(
      MyData[17]), .QN());
   DFFR_X1 \MyData_reg[16]  (.D(write_data[16]), .RN(n_1), .CK(n_0), .Q(
      MyData[16]), .QN());
   DFFR_X1 \MyData_reg[15]  (.D(write_data[15]), .RN(n_1), .CK(n_0), .Q(
      MyData[15]), .QN());
   DFFR_X1 \MyData_reg[14]  (.D(write_data[14]), .RN(n_1), .CK(n_0), .Q(
      MyData[14]), .QN());
   DFFR_X1 \MyData_reg[13]  (.D(write_data[13]), .RN(n_1), .CK(n_0), .Q(
      MyData[13]), .QN());
   DFFR_X1 \MyData_reg[12]  (.D(write_data[12]), .RN(n_1), .CK(n_0), .Q(
      MyData[12]), .QN());
   DFFR_X1 \MyData_reg[11]  (.D(write_data[11]), .RN(n_1), .CK(n_0), .Q(
      MyData[11]), .QN());
   DFFR_X1 \MyData_reg[10]  (.D(write_data[10]), .RN(n_1), .CK(n_0), .Q(
      MyData[10]), .QN());
   DFFR_X1 \MyData_reg[9]  (.D(write_data[9]), .RN(n_1), .CK(n_0), .Q(MyData[9]), 
      .QN());
   DFFR_X1 \MyData_reg[8]  (.D(write_data[8]), .RN(n_1), .CK(n_0), .Q(MyData[8]), 
      .QN());
   DFFR_X1 \MyData_reg[7]  (.D(write_data[7]), .RN(n_1), .CK(n_0), .Q(MyData[7]), 
      .QN());
   DFFR_X1 \MyData_reg[6]  (.D(write_data[6]), .RN(n_1), .CK(n_0), .Q(MyData[6]), 
      .QN());
   DFFR_X1 \MyData_reg[5]  (.D(write_data[5]), .RN(n_1), .CK(n_0), .Q(MyData[5]), 
      .QN());
   DFFR_X1 \MyData_reg[4]  (.D(write_data[4]), .RN(n_1), .CK(n_0), .Q(MyData[4]), 
      .QN());
   DFFR_X1 \MyData_reg[3]  (.D(write_data[3]), .RN(n_1), .CK(n_0), .Q(MyData[3]), 
      .QN());
   DFFR_X1 \MyData_reg[2]  (.D(write_data[2]), .RN(n_1), .CK(n_0), .Q(MyData[2]), 
      .QN());
   DFFR_X1 \MyData_reg[1]  (.D(write_data[1]), .RN(n_1), .CK(n_0), .Q(MyData[1]), 
      .QN());
   DFFR_X1 \MyData_reg[0]  (.D(write_data[0]), .RN(n_1), .CK(n_0), .Q(MyData[0]), 
      .QN());
endmodule

module AdderReg(i_Add1, i_Add2, result, write_enable, clk, rst);
   input [63:0]i_Add1;
   input [63:0]i_Add2;
   output [64:0]result;
   input write_enable;
   input clk;
   input rst;

   wire [64:0]Temp;

   ripple_adder adder (.i_add1(i_Add1), .i_add2(i_Add2), .o_result(Temp));
   Register RReg (.write_data(Temp), .write_enable(write_enable), .clk(clk), 
      .rst(rst), .MyData(result));
endmodule
