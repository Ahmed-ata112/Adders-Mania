/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Fri Nov  4 19:12:21 2022
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 272482328 */

/* blackbox module CLA_4bit_bbox */

/* blackbox module CLA_4bit_bbox_6 */

/* blackbox module CLA_4bit_bbox_5 */

/* blackbox module CLA_4bit_bbox_4 */

/* blackbox module CLA_4bit_bbox_3 */

/* blackbox module CLA_4bit_bbox_2 */

/* blackbox module CLA_4bit_bbox_1 */

/* blackbox module CLA_4bit_bbox_0 */

module CLA(in1, in2, cin, sum, cout, of);
   input [31:0]in1;
   input [31:0]in2;
   input cin;
   output [31:0]sum;
   output cout;
   output of;

   CLA_4bit_bbox cla1 (.a({in1[3], in1[2], in1[1], in1[0]}), .b({in2[3], in2[2], 
      in2[1], in2[0]}), .cin(1'b0), .sum({sum[3], sum[2], sum[1], sum[0]}), 
      .cout(n_0));
   CLA_4bit_bbox_6 cla2 (.a({in1[31], in1[31], in1[31], in1[31]}), .b({1'b0, 
      1'b0, 1'b0, 1'b0}), .cin(n_1), .sum({n_11, n_10, n_9, n_8}), .cout(n_7));
   CLA_4bit_bbox_5 genblk1_24_cla (.a({in1[31], in1[31], in1[31], in1[31]}), 
      .b({1'b0, 1'b0, 1'b0, 1'b0}), .cin(n_2), .sum({n_14, n_13, n_12, sum[24]}), 
      .cout(n_1));
   CLA_4bit_bbox_4 genblk1_20_cla (.a({in1[23], in1[22], in1[21], in1[20]}), 
      .b({in2[23], in2[22], in2[21], in2[20]}), .cin(n_3), .sum({sum[23], 
      sum[22], sum[21], sum[20]}), .cout(n_2));
   CLA_4bit_bbox_3 genblk1_16_cla (.a({in1[19], in1[18], in1[17], in1[16]}), 
      .b({in2[19], in2[18], in2[17], in2[16]}), .cin(n_4), .sum({sum[19], 
      sum[18], sum[17], sum[16]}), .cout(n_3));
   CLA_4bit_bbox_2 genblk1_12_cla (.a({in1[15], in1[14], in1[13], in1[12]}), 
      .b({in2[15], in2[14], in2[13], in2[12]}), .cin(n_5), .sum({sum[15], 
      sum[14], sum[13], sum[12]}), .cout(n_4));
   CLA_4bit_bbox_1 genblk1_8_cla (.a({in1[11], in1[10], in1[9], in1[8]}), 
      .b({in2[11], in2[10], in2[9], in2[8]}), .cin(n_6), .sum({sum[11], sum[10], 
      sum[9], sum[8]}), .cout(n_5));
   CLA_4bit_bbox_0 genblk1_4_cla (.a({in1[7], in1[6], in1[5], in1[4]}), .b({
      in2[7], in2[6], in2[5], in2[4]}), .cin(n_0), .sum({sum[7], sum[6], sum[5], 
      sum[4]}), .cout(n_6));
endmodule

module count_leading_zeros(valueIn, result);
   input [22:0]valueIn;
   output [4:0]result;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_22;
   wire n_0_27;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_28;
   wire n_0_29;

   AOI21_X1 i_0_0 (.A(valueIn[22]), .B1(n_0_40), .B2(n_0_0), .ZN(result[0]));
   OAI21_X1 i_0_1 (.A(n_0_39), .B1(valueIn[19]), .B2(n_0_1), .ZN(n_0_0));
   AOI21_X1 i_0_2 (.A(valueIn[18]), .B1(n_0_38), .B2(n_0_2), .ZN(n_0_1));
   OAI21_X1 i_0_3 (.A(n_0_37), .B1(valueIn[15]), .B2(n_0_3), .ZN(n_0_2));
   AOI21_X1 i_0_4 (.A(valueIn[14]), .B1(n_0_36), .B2(n_0_4), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(n_0_35), .B1(valueIn[11]), .B2(n_0_5), .ZN(n_0_4));
   AOI21_X1 i_0_6 (.A(valueIn[10]), .B1(n_0_34), .B2(n_0_6), .ZN(n_0_5));
   OAI21_X1 i_0_7 (.A(n_0_33), .B1(valueIn[7]), .B2(n_0_7), .ZN(n_0_6));
   AOI21_X1 i_0_8 (.A(valueIn[6]), .B1(n_0_32), .B2(n_0_8), .ZN(n_0_7));
   OAI21_X1 i_0_9 (.A(n_0_31), .B1(valueIn[3]), .B2(n_0_9), .ZN(n_0_8));
   AOI21_X1 i_0_10 (.A(valueIn[2]), .B1(n_0_30), .B2(valueIn[0]), .ZN(n_0_9));
   NOR3_X1 i_0_11 (.A1(valueIn[22]), .A2(valueIn[21]), .A3(n_0_10), .ZN(
      result[1]));
   NOR3_X1 i_0_12 (.A1(valueIn[20]), .A2(valueIn[19]), .A3(n_0_11), .ZN(n_0_10));
   NOR3_X1 i_0_13 (.A1(valueIn[18]), .A2(valueIn[17]), .A3(n_0_12), .ZN(n_0_11));
   NOR3_X1 i_0_14 (.A1(valueIn[16]), .A2(valueIn[15]), .A3(n_0_13), .ZN(n_0_12));
   NOR3_X1 i_0_15 (.A1(valueIn[14]), .A2(valueIn[13]), .A3(n_0_14), .ZN(n_0_13));
   AOI211_X1 i_0_16 (.A(valueIn[12]), .B(valueIn[11]), .C1(n_0_15), .C2(n_0_26), 
      .ZN(n_0_14));
   OAI21_X1 i_0_17 (.A(n_0_25), .B1(n_0_16), .B2(n_0_28), .ZN(n_0_15));
   NOR3_X1 i_0_18 (.A1(valueIn[4]), .A2(valueIn[3]), .A3(n_0_17), .ZN(n_0_16));
   NOR2_X1 i_0_19 (.A1(valueIn[2]), .A2(valueIn[1]), .ZN(n_0_17));
   AND3_X1 i_0_20 (.A1(n_0_22), .A2(n_0_24), .A3(n_0_23), .ZN(result[3]));
   NOR2_X1 i_0_21 (.A1(n_0_27), .A2(n_0_22), .ZN(result[4]));
   NAND3_X1 i_0_22 (.A1(n_0_29), .A2(n_0_26), .A3(n_0_25), .ZN(n_0_22));
   NAND2_X1 i_0_23 (.A1(n_0_23), .A2(n_0_24), .ZN(n_0_27));
   INV_X1 i_0_24 (.A(valueIn[1]), .ZN(n_0_30));
   INV_X1 i_0_25 (.A(valueIn[4]), .ZN(n_0_31));
   INV_X1 i_0_26 (.A(valueIn[5]), .ZN(n_0_32));
   INV_X1 i_0_27 (.A(valueIn[8]), .ZN(n_0_33));
   INV_X1 i_0_28 (.A(valueIn[9]), .ZN(n_0_34));
   INV_X1 i_0_29 (.A(valueIn[12]), .ZN(n_0_35));
   INV_X1 i_0_30 (.A(valueIn[13]), .ZN(n_0_36));
   INV_X1 i_0_31 (.A(valueIn[16]), .ZN(n_0_37));
   INV_X1 i_0_32 (.A(valueIn[17]), .ZN(n_0_38));
   INV_X1 i_0_33 (.A(valueIn[20]), .ZN(n_0_39));
   INV_X1 i_0_34 (.A(valueIn[21]), .ZN(n_0_40));
   AOI21_X1 i_0_35 (.A(n_0_21), .B1(n_0_24), .B2(n_0_18), .ZN(result[2]));
   OAI21_X1 i_0_36 (.A(n_0_29), .B1(n_0_20), .B2(n_0_19), .ZN(n_0_18));
   NAND2_X1 i_0_37 (.A1(n_0_26), .A2(n_0_25), .ZN(n_0_19));
   NOR3_X1 i_0_38 (.A1(valueIn[3]), .A2(n_0_28), .A3(valueIn[4]), .ZN(n_0_20));
   INV_X1 i_0_39 (.A(n_0_23), .ZN(n_0_21));
   NOR4_X1 i_0_40 (.A1(valueIn[22]), .A2(valueIn[21]), .A3(valueIn[20]), 
      .A4(valueIn[19]), .ZN(n_0_23));
   NOR4_X1 i_0_41 (.A1(valueIn[18]), .A2(valueIn[17]), .A3(valueIn[16]), 
      .A4(valueIn[15]), .ZN(n_0_24));
   NOR2_X1 i_0_42 (.A1(valueIn[8]), .A2(valueIn[7]), .ZN(n_0_25));
   NOR2_X1 i_0_43 (.A1(valueIn[10]), .A2(valueIn[9]), .ZN(n_0_26));
   OR2_X1 i_0_44 (.A1(valueIn[6]), .A2(valueIn[5]), .ZN(n_0_28));
   NOR4_X1 i_0_45 (.A1(valueIn[14]), .A2(valueIn[13]), .A3(valueIn[12]), 
      .A4(valueIn[11]), .ZN(n_0_29));
endmodule

module datapath__0_16(p_0, exp_Sum, p_1);
   output p_0;
   input [7:0]exp_Sum;
   input [21:0]p_1;

   NOR4_X1 i_0 (.A1(exp_Sum[7]), .A2(exp_Sum[6]), .A3(exp_Sum[5]), .A4(n_0), 
      .ZN(p_0));
   AOI21_X1 i_1 (.A(n_6), .B1(n_2), .B2(n_1), .ZN(n_0));
   AOI22_X1 i_2 (.A1(exp_Sum[4]), .A2(n_10), .B1(n_9), .B2(exp_Sum[3]), .ZN(n_1));
   OAI221_X1 i_3 (.A(n_3), .B1(n_8), .B2(exp_Sum[2]), .C1(exp_Sum[3]), .C2(n_9), 
      .ZN(n_2));
   NAND2_X1 i_4 (.A1(n_4), .A2(n_5), .ZN(n_3));
   AOI22_X1 i_5 (.A1(exp_Sum[2]), .A2(n_8), .B1(n_7), .B2(exp_Sum[1]), .ZN(n_4));
   OAI211_X1 i_6 (.A(exp_Sum[0]), .B(n_11), .C1(n_7), .C2(exp_Sum[1]), .ZN(n_5));
   NOR2_X1 i_7 (.A1(n_10), .A2(exp_Sum[4]), .ZN(n_6));
   INV_X1 i_8 (.A(p_1[1]), .ZN(n_7));
   INV_X1 i_9 (.A(p_1[2]), .ZN(n_8));
   INV_X1 i_10 (.A(p_1[3]), .ZN(n_9));
   INV_X1 i_11 (.A(p_1[4]), .ZN(n_10));
   INV_X1 i_12 (.A(p_1[11]), .ZN(n_11));
endmodule

module datapath__0_29(p_0, p_1);
   input [21:0]p_0;
   output [10:0]p_1;

   INV_X1 i_0 (.A(p_0[11]), .ZN(p_1[0]));
   HA_X1 i_1 (.A(p_0[1]), .B(p_0[11]), .CO(n_0), .S(p_1[1]));
   HA_X1 i_2 (.A(p_0[2]), .B(n_0), .CO(n_1), .S(p_1[2]));
   HA_X1 i_3 (.A(p_0[3]), .B(n_1), .CO(n_2), .S(p_1[3]));
   HA_X1 i_4 (.A(p_0[4]), .B(n_2), .CO(n_3), .S(p_1[4]));
endmodule

module datapath__0_34(mant_A, p_0);
   input [23:0]mant_A;
   output [31:0]p_0;

   XOR2_X1 i_0 (.A(mant_A[1]), .B(mant_A[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_21), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(mant_A[2]), .B1(mant_A[1]), .B2(mant_A[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(mant_A[3]), .B(n_21), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(mant_A[4]), .B(n_20), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(mant_A[5]), .B(n_19), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_18), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(mant_A[6]), .B1(n_19), .B2(mant_A[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(mant_A[7]), .B(n_18), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(mant_A[8]), .B(n_17), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_16), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(mant_A[9]), .B1(n_17), .B2(mant_A[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(mant_A[10]), .B(n_16), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(mant_A[11]), .B(n_15), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(mant_A[12]), .B(n_14), .Z(p_0[12]));
   XOR2_X1 i_15 (.A(mant_A[13]), .B(n_13), .Z(p_0[13]));
   XNOR2_X1 i_16 (.A(mant_A[14]), .B(n_12), .ZN(p_0[14]));
   XNOR2_X1 i_17 (.A(mant_A[15]), .B(n_11), .ZN(p_0[15]));
   XOR2_X1 i_18 (.A(mant_A[16]), .B(n_10), .Z(p_0[16]));
   XOR2_X1 i_19 (.A(mant_A[17]), .B(n_9), .Z(p_0[17]));
   XOR2_X1 i_20 (.A(mant_A[18]), .B(n_8), .Z(p_0[18]));
   AND2_X1 i_21 (.A1(n_7), .A2(n_3), .ZN(p_0[19]));
   OAI21_X1 i_22 (.A(mant_A[19]), .B1(n_8), .B2(mant_A[18]), .ZN(n_3));
   XOR2_X1 i_23 (.A(mant_A[20]), .B(n_7), .Z(p_0[20]));
   AND2_X1 i_24 (.A1(n_6), .A2(n_4), .ZN(p_0[21]));
   OAI21_X1 i_25 (.A(mant_A[21]), .B1(n_7), .B2(mant_A[20]), .ZN(n_4));
   XOR2_X1 i_26 (.A(mant_A[22]), .B(n_6), .Z(p_0[22]));
   AND2_X1 i_27 (.A1(p_0[31]), .A2(n_5), .ZN(p_0[23]));
   OAI21_X1 i_28 (.A(mant_A[23]), .B1(n_6), .B2(mant_A[22]), .ZN(n_5));
   OR3_X1 i_29 (.A1(n_6), .A2(mant_A[22]), .A3(mant_A[23]), .ZN(p_0[31]));
   OR3_X1 i_30 (.A1(n_7), .A2(mant_A[20]), .A3(mant_A[21]), .ZN(n_6));
   OR3_X1 i_31 (.A1(n_8), .A2(mant_A[18]), .A3(mant_A[19]), .ZN(n_7));
   OR2_X1 i_32 (.A1(n_9), .A2(mant_A[17]), .ZN(n_8));
   OR2_X1 i_33 (.A1(n_10), .A2(mant_A[16]), .ZN(n_9));
   NAND2_X1 i_34 (.A1(n_11), .A2(n_23), .ZN(n_10));
   NOR3_X1 i_35 (.A1(n_13), .A2(mant_A[13]), .A3(mant_A[14]), .ZN(n_11));
   NOR2_X1 i_36 (.A1(n_13), .A2(mant_A[13]), .ZN(n_12));
   OR2_X1 i_37 (.A1(n_14), .A2(mant_A[12]), .ZN(n_13));
   NAND2_X1 i_38 (.A1(n_15), .A2(n_22), .ZN(n_14));
   NOR2_X1 i_39 (.A1(n_16), .A2(mant_A[10]), .ZN(n_15));
   OR3_X1 i_40 (.A1(n_17), .A2(mant_A[8]), .A3(mant_A[9]), .ZN(n_16));
   OR2_X1 i_41 (.A1(n_18), .A2(mant_A[7]), .ZN(n_17));
   OR3_X1 i_42 (.A1(n_19), .A2(mant_A[5]), .A3(mant_A[6]), .ZN(n_18));
   OR2_X1 i_43 (.A1(n_20), .A2(mant_A[4]), .ZN(n_19));
   OR2_X1 i_44 (.A1(n_21), .A2(mant_A[3]), .ZN(n_20));
   OR3_X1 i_45 (.A1(mant_A[2]), .A2(mant_A[1]), .A3(mant_A[0]), .ZN(n_21));
   INV_X1 i_46 (.A(mant_A[11]), .ZN(n_22));
   INV_X1 i_47 (.A(mant_A[15]), .ZN(n_23));
endmodule

module fp_adder(A, B, Sum, overflow, underflow);
   input [31:0]A;
   input [31:0]B;
   output [31:0]Sum;
   output overflow;
   output underflow;

   wire [4:0]num_leading_zeros;
   wire n_0_5;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_0_7;
   wire n_0_0_0;
   wire n_0_0_8;
   wire n_0_0_1;
   wire n_0_0_9;
   wire n_0_0_2;
   wire n_0_0_10;
   wire n_0_0_3;
   wire n_0_0_11;
   wire n_0_0_4;
   wire n_0_0_12;
   wire n_0_0_5;
   wire n_0_0_13;
   wire n_0_0_6;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_127;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire [31:0]mant_A;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_231;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_0_246;
   wire n_0_0_247;
   wire n_0_0_248;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_0_253;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_0_260;
   wire n_0_0_261;
   wire [7:0]exp_Sum;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_30;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_31;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_32;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_0_288;
   wire n_0_0_289;
   wire n_0_33;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_0_294;
   wire n_0_34;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_35;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_0_304;
   wire n_0_0_305;
   wire n_0_37;
   wire n_0_0_311;
   wire n_0_38;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_39;
   wire n_0_0_320;
   wire n_0_0_321;
   wire n_0_0_322;
   wire n_0_40;
   wire n_0_0_328;
   wire n_0_0_329;
   wire n_0_0_330;
   wire n_0_0_331;
   wire n_0_0_332;
   wire n_0_41;
   wire n_0_0_334;
   wire n_0_0_335;
   wire n_0_0_336;
   wire n_0_42;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_341;
   wire n_0_43;
   wire n_0_0_342;
   wire n_0_0_343;
   wire n_0_0_344;
   wire n_0_44;
   wire n_0_0_346;
   wire n_0_0_347;
   wire n_0_0_348;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_351;
   wire n_0_0_355;
   wire n_0_45;
   wire n_0_0_356;
   wire n_0_0_357;
   wire n_0_0_358;
   wire n_0_46;
   wire n_0_0_359;
   wire n_0_0_360;
   wire n_0_47;
   wire n_0_0_363;
   wire n_0_0_364;
   wire n_0_0_365;
   wire n_0_48;
   wire n_0_0_367;
   wire n_0_0_368;
   wire n_0_0_370;
   wire n_0_0_371;
   wire n_0_0_372;
   wire n_0_0_373;
   wire n_0_49;
   wire n_0_0_376;
   wire n_0_0_377;
   wire n_0_0_378;
   wire n_0_50;
   wire n_0_0_379;
   wire n_0_0_380;
   wire n_0_51;
   wire n_0_0_381;
   wire n_0_0_382;
   wire n_0_0_396;
   wire n_0_0_397;
   wire n_0_0_398;
   wire n_0_0_399;
   wire n_0_0_400;
   wire n_0_0_401;
   wire n_0_0_402;
   wire n_0_0_403;
   wire n_0_0_404;
   wire n_0_0_405;
   wire n_0_0_406;
   wire n_0_0_407;
   wire n_0_0_408;
   wire n_0_0_409;
   wire n_0_0_410;
   wire n_0_0_411;
   wire n_0_0_412;
   wire n_0_0_413;
   wire n_0_0_414;
   wire n_0_0_415;
   wire n_0_0_416;
   wire n_0_0_417;
   wire n_0_0_418;
   wire n_0_0_419;
   wire n_0_0_420;
   wire n_0_0_426;
   wire n_0_0_431;
   wire n_0_0_432;
   wire n_0_0_437;
   wire n_0_0_438;
   wire n_0_0_443;
   wire n_0_0_444;
   wire n_0_0_445;
   wire n_0_0_446;
   wire n_0_0_447;
   wire n_0_0_448;
   wire n_0_0_449;
   wire n_0_0_451;
   wire n_0_0_452;
   wire n_0_0_453;
   wire n_0_0_454;
   wire n_0_0_455;
   wire n_0_0_456;
   wire n_0_0_457;
   wire n_0_0_458;
   wire n_0_0_459;
   wire n_0_0_460;
   wire n_0_0_461;
   wire n_0_0_462;
   wire n_0_0_463;
   wire n_0_0_464;
   wire n_0_0_465;
   wire n_0_0_466;
   wire n_0_0_467;
   wire n_0_0_468;
   wire n_0_0_469;
   wire n_0_0_472;
   wire n_0_0_473;
   wire n_0_0_474;
   wire n_0_0_475;
   wire n_0_0_476;
   wire n_0_0_477;
   wire n_0_0_478;
   wire n_0_0_479;
   wire n_0_0_480;
   wire n_0_0_481;
   wire n_0_0_482;
   wire n_0_0_483;
   wire n_0_0_485;
   wire n_0_0_486;
   wire n_0_0_487;
   wire n_0_0_488;
   wire n_0_0_489;
   wire n_0_0_490;
   wire n_0_0_491;
   wire n_0_0_494;
   wire n_0_0_496;
   wire n_0_0_497;
   wire n_0_0_498;
   wire n_0_0_499;
   wire n_0_0_500;
   wire n_0_0_501;
   wire n_0_0_502;
   wire n_0_0_504;
   wire n_0_0_515;
   wire n_0_0_95;
   wire n_0_0_532;
   wire n_0_0_563;
   wire n_0_0_564;
   wire n_0_0_578;
   wire n_0_0_579;
   wire n_0_0_580;
   wire n_0_0_581;
   wire n_0_0_582;
   wire n_0_0_583;
   wire n_0_0_584;
   wire n_0_0_585;
   wire n_0_0_586;
   wire n_0_0_587;
   wire n_0_0_588;
   wire n_0_0_96;
   wire n_0_0_603;
   wire n_0_0_604;
   wire n_0_0_605;
   wire n_0_0_606;
   wire n_0_0_607;
   wire n_0_0_608;
   wire n_0_0_609;
   wire n_0_0_610;
   wire n_0_0_611;
   wire n_0_0_612;
   wire n_0_0_613;
   wire n_0_0_99;
   wire n_0_0_94;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_0_312;
   wire n_0_0_313;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_0_319;
   wire n_0_0_323;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_333;
   wire n_0_0_345;
   wire n_0_0_352;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_0_361;
   wire n_0_0_362;
   wire n_0_36;
   wire n_0_0_366;
   wire n_0_0_369;
   wire n_0_0_374;
   wire n_0_0_375;
   wire n_0_0_383;
   wire n_0_0_384;
   wire n_0_0_385;
   wire n_0_0_386;
   wire n_0_0_387;
   wire n_0_0_388;
   wire n_0_0_389;
   wire n_0_0_390;
   wire n_0_0_391;
   wire n_0_0_392;
   wire n_0_0_393;
   wire n_0_0_394;
   wire n_0_0_395;
   wire n_0_0_421;
   wire n_0_0_422;
   wire n_0_0_423;
   wire n_0_0_424;
   wire n_0_0_425;
   wire n_0_0_427;
   wire n_0_0_428;
   wire n_0_0_429;
   wire n_0_0_430;
   wire n_0_0_433;
   wire n_0_0_434;
   wire n_0_0_435;
   wire n_0_0_436;
   wire n_0_0_439;
   wire n_0_0_440;
   wire n_0_0_441;
   wire n_0_0_442;
   wire n_0_0_450;
   wire n_0_0_470;
   wire n_0_0_471;
   wire n_0_0_484;
   wire n_0_0_492;
   wire n_0_0_493;
   wire n_0_0_495;
   wire n_0_0_503;
   wire n_0_0_505;
   wire n_0_0_506;
   wire n_0_0_507;
   wire n_0_0_508;
   wire n_0_0_509;
   wire n_0_0_510;
   wire n_0_0_511;
   wire n_0_0_512;
   wire n_0_0_513;
   wire n_0_0_514;
   wire n_0_0_516;
   wire n_0_52;
   wire n_0_0_517;
   wire n_0_0_518;
   wire n_0_0_519;
   wire n_0_0_520;
   wire n_0_0_521;
   wire n_0_0_522;
   wire n_0_0_523;
   wire n_0_0_524;
   wire n_0_0_525;
   wire n_0_0_526;
   wire n_0_0_527;
   wire n_0_0_528;
   wire n_0_0_529;
   wire n_0_0_530;
   wire n_0_0_531;
   wire n_0_0_533;
   wire n_0_0_534;
   wire n_0_0_535;
   wire n_0_0_536;
   wire n_0_0_537;
   wire n_0_0_538;
   wire n_0_0_539;
   wire n_0_0_540;
   wire n_0_0_541;
   wire n_0_0_542;
   wire n_0_0_543;
   wire n_0_0_544;
   wire n_0_0_545;
   wire n_0_0_546;
   wire n_0_0_547;
   wire n_0_0_548;
   wire n_0_0_549;
   wire n_0_0_550;
   wire n_0_0_551;
   wire n_0_0_552;
   wire n_0_0_553;
   wire n_0_0_554;
   wire n_0_0_555;
   wire n_0_0_556;
   wire n_0_0_557;
   wire n_0_0_558;
   wire n_0_0_559;
   wire n_0_0_560;
   wire n_0_0_561;
   wire n_0_0_562;
   wire n_0_0_565;
   wire n_0_0_566;
   wire n_0_0_567;
   wire n_0_0_568;
   wire n_0_0_569;
   wire n_0_0_570;
   wire n_0_0_571;
   wire n_0_0_572;
   wire n_0_0_573;
   wire n_0_0_574;
   wire n_0_0_575;
   wire n_0_0_576;
   wire n_0_0_577;
   wire n_0_0_589;
   wire n_0_0_590;
   wire n_0_0_591;
   wire n_0_0_592;
   wire n_0_0_593;
   wire n_0_0_594;
   wire n_0_0_595;
   wire n_0_0_596;
   wire n_0_0_597;
   wire n_0_0_598;
   wire n_0_0_599;
   wire n_0_0_600;
   wire n_0_0_601;
   wire n_0_0_602;
   wire n_0_0_614;
   wire n_0_0_615;
   wire n_0_0_616;
   wire n_0_0_617;

   CLA CLA_dut (.in1({mant_A[31], uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, 
      mant_A[23], mant_A[22], mant_A[21], mant_A[20], mant_A[19], mant_A[18], 
      mant_A[17], mant_A[16], mant_A[15], mant_A[14], mant_A[13], mant_A[12], 
      mant_A[11], mant_A[10], mant_A[9], mant_A[8], mant_A[7], mant_A[6], 
      mant_A[5], mant_A[4], mant_A[3], mant_A[2], mant_A[1], mant_A[0]}), 
      .in2({uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, n_48, n_46, 
      n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, n_36, n_35, n_34, 
      n_33, n_32, n_31, n_30, n_47, n_29, n_28, n_27, n_26, n_25}), .cin(), 
      .sum({uc_15, uc_16, uc_17, uc_18, uc_19, uc_20, uc_21, n_24, n_23, n_22, 
      n_21, n_20, n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, 
      n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, n_1, n_0}), .cout(), .of());
   count_leading_zeros count_leading_zeros_instance (.valueIn({n_22, n_21, n_20, 
      n_19, n_18, n_17, n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, 
      n_6, n_5, n_4, n_3, n_2, n_1, n_0}), .result(num_leading_zeros));
   datapath__0_16 i_0_5 (.p_0(n_0_5), .exp_Sum(exp_Sum), .p_1({1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, num_leading_zeros[0], 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, num_leading_zeros[4], num_leading_zeros[3], 
      num_leading_zeros[2], num_leading_zeros[1], 1'b1}));
   datapath__0_29 i_0_17 (.p_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, num_leading_zeros[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      num_leading_zeros[4], num_leading_zeros[3], num_leading_zeros[2], 
      num_leading_zeros[1], 1'b1}), .p_1({uc_22, uc_23, uc_24, uc_25, uc_26, 
      uc_27, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0}));
   datapath__0_34 i_0_22 (.mant_A({n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, 
      n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, 
      n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, n_0_30, 
      mant_A[0]}), .p_0({n_0_29, uc_28, uc_29, uc_30, uc_31, uc_32, uc_33, uc_34, 
      n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, 
      n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, 
      n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, uc_35}));
   HA_X1 i_0_0_0 (.A(n_24), .B(exp_Sum[0]), .CO(n_0_0_0), .S(n_0_0_7));
   HA_X1 i_0_0_1 (.A(exp_Sum[1]), .B(n_0_0_0), .CO(n_0_0_1), .S(n_0_0_8));
   HA_X1 i_0_0_2 (.A(exp_Sum[2]), .B(n_0_0_1), .CO(n_0_0_2), .S(n_0_0_9));
   HA_X1 i_0_0_3 (.A(exp_Sum[3]), .B(n_0_0_2), .CO(n_0_0_3), .S(n_0_0_10));
   HA_X1 i_0_0_4 (.A(exp_Sum[4]), .B(n_0_0_3), .CO(n_0_0_4), .S(n_0_0_11));
   HA_X1 i_0_0_5 (.A(exp_Sum[5]), .B(n_0_0_4), .CO(n_0_0_5), .S(n_0_0_12));
   HA_X1 i_0_0_6 (.A(exp_Sum[6]), .B(n_0_0_5), .CO(n_0_0_6), .S(n_0_0_13));
   INV_X1 i_0_0_7 (.A(n_0_0_14), .ZN(Sum[0]));
   AOI22_X1 i_0_0_8 (.A1(n_0), .A2(n_0_0_17), .B1(n_1), .B2(n_0_0_136), .ZN(
      n_0_0_14));
   OAI21_X1 i_0_0_9 (.A(n_0_0_15), .B1(n_0_0_134), .B2(n_0_0_16), .ZN(Sum[1]));
   AOI22_X1 i_0_0_10 (.A1(n_1), .A2(n_0_0_17), .B1(n_2), .B2(n_0_0_136), 
      .ZN(n_0_0_15));
   NAND2_X1 i_0_0_11 (.A1(n_0), .A2(n_0_0_25), .ZN(n_0_0_16));
   INV_X1 i_0_0_12 (.A(n_0_0_18), .ZN(n_0_0_17));
   AOI21_X1 i_0_0_13 (.A(n_0_0_137), .B1(n_0_0_116), .B2(n_0_0_25), .ZN(n_0_0_18));
   OAI221_X1 i_0_0_14 (.A(n_0_0_19), .B1(n_0_0_134), .B2(n_0_0_20), .C1(
      n_0_0_115), .C2(n_0_0_21), .ZN(Sum[2]));
   AOI22_X1 i_0_0_15 (.A1(n_3), .A2(n_0_0_136), .B1(n_2), .B2(n_0_0_137), 
      .ZN(n_0_0_19));
   NAND2_X1 i_0_0_16 (.A1(n_1), .A2(n_0_0_25), .ZN(n_0_0_20));
   OAI221_X1 i_0_0_17 (.A(n_0_0_22), .B1(n_0_0_134), .B2(n_0_0_21), .C1(
      n_0_0_115), .C2(n_0_0_24), .ZN(Sum[3]));
   AOI22_X1 i_0_0_18 (.A1(n_0), .A2(n_0_0_34), .B1(n_2), .B2(n_0_0_25), .ZN(
      n_0_0_21));
   AOI22_X1 i_0_0_19 (.A1(n_3), .A2(n_0_0_137), .B1(n_4), .B2(n_0_0_136), 
      .ZN(n_0_0_22));
   OAI21_X1 i_0_0_20 (.A(n_0_0_23), .B1(n_0_0_134), .B2(n_0_0_24), .ZN(Sum[4]));
   AOI222_X1 i_0_0_21 (.A1(n_5), .A2(n_0_0_136), .B1(n_4), .B2(n_0_0_137), 
      .C1(n_0_0_116), .C2(n_0_0_27), .ZN(n_0_0_23));
   AOI22_X1 i_0_0_22 (.A1(n_1), .A2(n_0_0_34), .B1(n_3), .B2(n_0_0_25), .ZN(
      n_0_0_24));
   AND2_X1 i_0_0_23 (.A1(n_0_0_125), .A2(n_0_0_113), .ZN(n_0_0_25));
   NAND2_X1 i_0_0_24 (.A1(n_0_0_29), .A2(n_0_0_26), .ZN(Sum[5]));
   AOI22_X1 i_0_0_25 (.A1(n_0_0_133), .A2(n_0_0_27), .B1(n_5), .B2(n_0_0_137), 
      .ZN(n_0_0_26));
   OAI21_X1 i_0_0_26 (.A(n_0_0_28), .B1(n_0_1), .B2(n_0_0_37), .ZN(n_0_0_27));
   NAND2_X1 i_0_0_27 (.A1(n_2), .A2(n_0_0_34), .ZN(n_0_0_28));
   AOI22_X1 i_0_0_28 (.A1(n_6), .A2(n_0_0_136), .B1(n_0_0_116), .B2(n_0_0_32), 
      .ZN(n_0_0_29));
   NAND2_X1 i_0_0_29 (.A1(n_0_0_31), .A2(n_0_0_30), .ZN(Sum[6]));
   AOI22_X1 i_0_0_30 (.A1(n_6), .A2(n_0_0_137), .B1(n_0_0_116), .B2(n_0_0_36), 
      .ZN(n_0_0_30));
   AOI22_X1 i_0_0_31 (.A1(n_0_0_133), .A2(n_0_0_32), .B1(n_7), .B2(n_0_0_136), 
      .ZN(n_0_0_31));
   OAI21_X1 i_0_0_32 (.A(n_0_0_33), .B1(n_0_1), .B2(n_0_0_41), .ZN(n_0_0_32));
   NAND2_X1 i_0_0_33 (.A1(n_3), .A2(n_0_0_34), .ZN(n_0_0_33));
   AND2_X1 i_0_0_34 (.A1(n_0_1), .A2(n_0_0_113), .ZN(n_0_0_34));
   NAND2_X1 i_0_0_35 (.A1(n_0_0_38), .A2(n_0_0_35), .ZN(Sum[7]));
   AOI22_X1 i_0_0_36 (.A1(n_0_0_133), .A2(n_0_0_36), .B1(n_7), .B2(n_0_0_137), 
      .ZN(n_0_0_35));
   OAI22_X1 i_0_0_37 (.A1(n_0_1), .A2(n_0_0_46), .B1(n_0_0_125), .B2(n_0_0_37), 
      .ZN(n_0_0_36));
   AOI22_X1 i_0_0_38 (.A1(n_4), .A2(n_0_0_113), .B1(n_0), .B2(n_0_0_87), 
      .ZN(n_0_0_37));
   AOI22_X1 i_0_0_39 (.A1(n_8), .A2(n_0_0_136), .B1(n_0_0_116), .B2(n_0_0_40), 
      .ZN(n_0_0_38));
   NAND2_X1 i_0_0_40 (.A1(n_0_0_42), .A2(n_0_0_39), .ZN(Sum[8]));
   AOI22_X1 i_0_0_41 (.A1(n_0_0_116), .A2(n_0_0_45), .B1(n_0_0_133), .B2(
      n_0_0_40), .ZN(n_0_0_39));
   OAI22_X1 i_0_0_42 (.A1(n_0_1), .A2(n_0_0_49), .B1(n_0_0_125), .B2(n_0_0_41), 
      .ZN(n_0_0_40));
   AOI22_X1 i_0_0_43 (.A1(n_5), .A2(n_0_0_113), .B1(n_1), .B2(n_0_0_87), 
      .ZN(n_0_0_41));
   AOI22_X1 i_0_0_44 (.A1(n_9), .A2(n_0_0_136), .B1(n_8), .B2(n_0_0_137), 
      .ZN(n_0_0_42));
   NAND2_X1 i_0_0_45 (.A1(n_0_0_44), .A2(n_0_0_43), .ZN(Sum[9]));
   AOI22_X1 i_0_0_46 (.A1(n_9), .A2(n_0_0_137), .B1(n_0_0_116), .B2(n_0_0_48), 
      .ZN(n_0_0_43));
   AOI22_X1 i_0_0_47 (.A1(n_0_0_133), .A2(n_0_0_45), .B1(n_10), .B2(n_0_0_136), 
      .ZN(n_0_0_44));
   OAI22_X1 i_0_0_48 (.A1(n_0_1), .A2(n_0_0_53), .B1(n_0_0_125), .B2(n_0_0_46), 
      .ZN(n_0_0_45));
   AOI22_X1 i_0_0_49 (.A1(n_6), .A2(n_0_0_113), .B1(n_2), .B2(n_0_0_87), 
      .ZN(n_0_0_46));
   NAND2_X1 i_0_0_50 (.A1(n_0_0_50), .A2(n_0_0_47), .ZN(Sum[10]));
   AOI22_X1 i_0_0_51 (.A1(n_10), .A2(n_0_0_137), .B1(n_0_0_133), .B2(n_0_0_48), 
      .ZN(n_0_0_47));
   OAI22_X1 i_0_0_52 (.A1(n_0_0_125), .A2(n_0_0_49), .B1(n_0_1), .B2(n_0_0_58), 
      .ZN(n_0_0_48));
   AOI22_X1 i_0_0_53 (.A1(n_7), .A2(n_0_0_113), .B1(n_3), .B2(n_0_0_87), 
      .ZN(n_0_0_49));
   AOI22_X1 i_0_0_54 (.A1(n_0_0_116), .A2(n_0_0_52), .B1(n_11), .B2(n_0_0_136), 
      .ZN(n_0_0_50));
   NAND2_X1 i_0_0_55 (.A1(n_0_0_54), .A2(n_0_0_51), .ZN(Sum[11]));
   AOI22_X1 i_0_0_56 (.A1(n_0_0_133), .A2(n_0_0_52), .B1(n_0_0_116), .B2(
      n_0_0_57), .ZN(n_0_0_51));
   OAI22_X1 i_0_0_57 (.A1(n_0_1), .A2(n_0_0_62), .B1(n_0_0_125), .B2(n_0_0_53), 
      .ZN(n_0_0_52));
   AOI222_X1 i_0_0_58 (.A1(n_8), .A2(n_0_0_113), .B1(n_0), .B2(n_0_0_119), 
      .C1(n_4), .C2(n_0_0_87), .ZN(n_0_0_53));
   AOI22_X1 i_0_0_59 (.A1(n_11), .A2(n_0_0_137), .B1(n_12), .B2(n_0_0_136), 
      .ZN(n_0_0_54));
   NAND2_X1 i_0_0_60 (.A1(n_0_0_56), .A2(n_0_0_55), .ZN(Sum[12]));
   AOI22_X1 i_0_0_61 (.A1(n_12), .A2(n_0_0_137), .B1(n_0_0_116), .B2(n_0_0_60), 
      .ZN(n_0_0_55));
   AOI22_X1 i_0_0_62 (.A1(n_0_0_133), .A2(n_0_0_57), .B1(n_13), .B2(n_0_0_136), 
      .ZN(n_0_0_56));
   OAI22_X1 i_0_0_63 (.A1(n_0_1), .A2(n_0_0_68), .B1(n_0_0_125), .B2(n_0_0_58), 
      .ZN(n_0_0_57));
   AOI222_X1 i_0_0_64 (.A1(n_9), .A2(n_0_0_113), .B1(n_1), .B2(n_0_0_119), 
      .C1(n_5), .C2(n_0_0_87), .ZN(n_0_0_58));
   NAND2_X1 i_0_0_65 (.A1(n_0_0_63), .A2(n_0_0_59), .ZN(Sum[13]));
   AOI22_X1 i_0_0_66 (.A1(n_13), .A2(n_0_0_137), .B1(n_0_0_133), .B2(n_0_0_60), 
      .ZN(n_0_0_59));
   OAI21_X1 i_0_0_67 (.A(n_0_0_61), .B1(n_0_0_125), .B2(n_0_0_62), .ZN(n_0_0_60));
   NAND2_X1 i_0_0_68 (.A1(n_0_0_125), .A2(n_0_0_71), .ZN(n_0_0_61));
   AOI222_X1 i_0_0_69 (.A1(n_10), .A2(n_0_0_113), .B1(n_2), .B2(n_0_0_119), 
      .C1(n_6), .C2(n_0_0_87), .ZN(n_0_0_62));
   AOI22_X1 i_0_0_70 (.A1(n_0_0_116), .A2(n_0_0_66), .B1(n_14), .B2(n_0_0_136), 
      .ZN(n_0_0_63));
   OAI211_X1 i_0_0_71 (.A(n_0_0_64), .B(n_0_0_65), .C1(n_0_0_115), .C2(n_0_0_70), 
      .ZN(Sum[14]));
   NAND2_X1 i_0_0_72 (.A1(n_14), .A2(n_0_0_137), .ZN(n_0_0_64));
   AOI22_X1 i_0_0_73 (.A1(n_15), .A2(n_0_0_136), .B1(n_0_0_133), .B2(n_0_0_66), 
      .ZN(n_0_0_65));
   OAI21_X1 i_0_0_74 (.A(n_0_0_67), .B1(n_0_0_125), .B2(n_0_0_68), .ZN(n_0_0_66));
   NAND2_X1 i_0_0_75 (.A1(n_0_0_125), .A2(n_0_0_77), .ZN(n_0_0_67));
   AOI222_X1 i_0_0_76 (.A1(n_11), .A2(n_0_0_113), .B1(n_3), .B2(n_0_0_119), 
      .C1(n_7), .C2(n_0_0_87), .ZN(n_0_0_68));
   OAI221_X1 i_0_0_77 (.A(n_0_0_69), .B1(n_0_0_134), .B2(n_0_0_70), .C1(
      n_0_0_115), .C2(n_0_0_76), .ZN(Sum[15]));
   AOI22_X1 i_0_0_78 (.A1(n_16), .A2(n_0_0_136), .B1(n_15), .B2(n_0_0_137), 
      .ZN(n_0_0_69));
   AOI22_X1 i_0_0_79 (.A1(n_0_0_125), .A2(n_0_0_80), .B1(n_0_1), .B2(n_0_0_71), 
      .ZN(n_0_0_70));
   OAI21_X1 i_0_0_80 (.A(n_0_0_72), .B1(n_0_2), .B2(n_0_0_92), .ZN(n_0_0_71));
   AOI22_X1 i_0_0_81 (.A1(n_0), .A2(n_0_0_86), .B1(n_8), .B2(n_0_0_87), .ZN(
      n_0_0_72));
   OAI211_X1 i_0_0_82 (.A(n_0_0_74), .B(n_0_0_73), .C1(n_0_0_115), .C2(n_0_0_79), 
      .ZN(Sum[16]));
   NAND2_X1 i_0_0_83 (.A1(n_16), .A2(n_0_0_137), .ZN(n_0_0_73));
   AOI22_X1 i_0_0_84 (.A1(n_0_0_133), .A2(n_0_0_75), .B1(n_17), .B2(n_0_0_136), 
      .ZN(n_0_0_74));
   INV_X1 i_0_0_85 (.A(n_0_0_76), .ZN(n_0_0_75));
   AOI22_X1 i_0_0_86 (.A1(n_0_0_125), .A2(n_0_0_84), .B1(n_0_1), .B2(n_0_0_77), 
      .ZN(n_0_0_76));
   OAI21_X1 i_0_0_87 (.A(n_0_0_78), .B1(n_0_2), .B2(n_0_0_109), .ZN(n_0_0_77));
   AOI22_X1 i_0_0_88 (.A1(n_1), .A2(n_0_0_86), .B1(n_9), .B2(n_0_0_87), .ZN(
      n_0_0_78));
   OAI221_X1 i_0_0_89 (.A(n_0_0_82), .B1(n_0_0_134), .B2(n_0_0_79), .C1(
      n_0_0_115), .C2(n_0_0_83), .ZN(Sum[17]));
   AOI22_X1 i_0_0_90 (.A1(n_0_0_125), .A2(n_0_0_91), .B1(n_0_1), .B2(n_0_0_80), 
      .ZN(n_0_0_79));
   OAI21_X1 i_0_0_91 (.A(n_0_0_81), .B1(n_0_2), .B2(n_0_0_196), .ZN(n_0_0_80));
   AOI22_X1 i_0_0_92 (.A1(n_10), .A2(n_0_0_87), .B1(n_2), .B2(n_0_0_86), 
      .ZN(n_0_0_81));
   AOI22_X1 i_0_0_93 (.A1(n_17), .A2(n_0_0_137), .B1(n_18), .B2(n_0_0_136), 
      .ZN(n_0_0_82));
   OAI221_X1 i_0_0_94 (.A(n_0_0_88), .B1(n_0_0_115), .B2(n_0_0_90), .C1(
      n_0_0_134), .C2(n_0_0_83), .ZN(Sum[18]));
   AOI22_X1 i_0_0_95 (.A1(n_0_1), .A2(n_0_0_84), .B1(n_0_0_125), .B2(n_0_0_101), 
      .ZN(n_0_0_83));
   OAI21_X1 i_0_0_96 (.A(n_0_0_85), .B1(n_0_2), .B2(n_0_0_112), .ZN(n_0_0_84));
   AOI22_X1 i_0_0_97 (.A1(n_11), .A2(n_0_0_87), .B1(n_3), .B2(n_0_0_86), 
      .ZN(n_0_0_85));
   NOR3_X1 i_0_0_98 (.A1(n_0_4), .A2(n_0_0_128), .A3(n_0_0_126), .ZN(n_0_0_86));
   NOR3_X1 i_0_0_99 (.A1(n_0_4), .A2(n_0_3), .A3(n_0_0_126), .ZN(n_0_0_87));
   AOI22_X1 i_0_0_100 (.A1(n_19), .A2(n_0_0_136), .B1(n_18), .B2(n_0_0_137), 
      .ZN(n_0_0_88));
   OAI221_X1 i_0_0_101 (.A(n_0_0_89), .B1(n_0_0_134), .B2(n_0_0_90), .C1(
      n_0_0_115), .C2(n_0_0_100), .ZN(Sum[19]));
   AOI22_X1 i_0_0_102 (.A1(n_20), .A2(n_0_0_136), .B1(n_19), .B2(n_0_0_137), 
      .ZN(n_0_0_89));
   AOI22_X1 i_0_0_103 (.A1(n_0_0_125), .A2(n_0_0_195), .B1(n_0_1), .B2(n_0_0_91), 
      .ZN(n_0_0_90));
   OAI22_X1 i_0_0_104 (.A1(n_0_2), .A2(n_0_0_194), .B1(n_0_0_126), .B2(n_0_0_92), 
      .ZN(n_0_0_91));
   AOI22_X1 i_0_0_105 (.A1(n_4), .A2(n_0_0_120), .B1(n_12), .B2(n_0_0_114), 
      .ZN(n_0_0_92));
   OAI211_X1 i_0_0_106 (.A(n_0_0_97), .B(n_0_0_93), .C1(n_0_0_134), .C2(
      n_0_0_100), .ZN(Sum[20]));
   AOI22_X1 i_0_0_107 (.A1(n_20), .A2(n_0_0_137), .B1(n_0_0_116), .B2(n_0_0_130), 
      .ZN(n_0_0_93));
   NAND2_X1 i_0_0_108 (.A1(n_21), .A2(n_0_0_136), .ZN(n_0_0_97));
   NAND2_X1 i_0_0_109 (.A1(n_0_0_103), .A2(n_0_0_98), .ZN(Sum[21]));
   AOI22_X1 i_0_0_110 (.A1(n_0_0_133), .A2(n_0_0_130), .B1(n_21), .B2(n_0_0_137), 
      .ZN(n_0_0_98));
   AOI22_X1 i_0_0_111 (.A1(n_22), .A2(n_0_0_136), .B1(n_0_0_117), .B2(n_0_0_116), 
      .ZN(n_0_0_103));
   NAND2_X1 i_0_0_112 (.A1(n_0_0_135), .A2(n_0_0_104), .ZN(Sum[22]));
   AOI21_X1 i_0_0_113 (.A(n_0_0_105), .B1(n_0_0_133), .B2(n_0_0_117), .ZN(
      n_0_0_104));
   AOI221_X1 i_0_0_114 (.A(n_0_0_115), .B1(n_0_0_125), .B2(n_0_0_106), .C1(n_0_1), 
      .C2(n_0_0_132), .ZN(n_0_0_105));
   AOI21_X1 i_0_0_115 (.A(n_0_0_107), .B1(n_22), .B2(n_0_0_113), .ZN(n_0_0_106));
   OAI21_X1 i_0_0_116 (.A(n_0_0_108), .B1(n_0_0_126), .B2(n_0_0_197), .ZN(
      n_0_0_107));
   AOI22_X1 i_0_0_117 (.A1(n_14), .A2(n_0_0_119), .B1(n_6), .B2(n_0_0_121), 
      .ZN(n_0_0_108));
   INV_X1 i_0_0_118 (.A(n_0_0_116), .ZN(n_0_0_115));
   NOR2_X1 i_0_0_119 (.A1(n_0_0), .A2(n_0_0_228), .ZN(n_0_0_116));
   INV_X1 i_0_0_120 (.A(n_0_0_118), .ZN(n_0_0_117));
   OAI22_X1 i_0_0_121 (.A1(n_0_0_125), .A2(n_0_0_110), .B1(n_0_1), .B2(n_0_0_123), 
      .ZN(n_0_0_118));
   OAI211_X1 i_0_0_122 (.A(n_0_0_127), .B(n_0_0_124), .C1(n_0_0_126), .C2(
      n_0_0_102), .ZN(n_0_0_123));
   AOI22_X1 i_0_0_123 (.A1(n_21), .A2(n_0_0_113), .B1(n_5), .B2(n_0_0_121), 
      .ZN(n_0_0_124));
   NAND2_X1 i_0_0_124 (.A1(n_13), .A2(n_0_0_119), .ZN(n_0_0_127));
   INV_X1 i_0_0_125 (.A(n_0_0_134), .ZN(n_0_0_133));
   NAND2_X1 i_0_0_126 (.A1(n_0_0), .A2(n_0_0_229), .ZN(n_0_0_134));
   AOI22_X1 i_0_0_127 (.A1(n_22), .A2(n_0_0_137), .B1(n_23), .B2(n_0_0_136), 
      .ZN(n_0_0_135));
   AND3_X1 i_0_0_128 (.A1(n_24), .A2(n_0_0_232), .A3(n_0_0_225), .ZN(n_0_0_136));
   OAI21_X1 i_0_0_129 (.A(n_0_0_154), .B1(n_24), .B2(n_0_0_233), .ZN(n_0_0_137));
   INV_X1 i_0_0_130 (.A(n_0_0_138), .ZN(Sum[23]));
   AOI222_X1 i_0_0_131 (.A1(n_0_0_7), .A2(n_0_0_232), .B1(exp_Sum[0]), .B2(
      n_0_0_153), .C1(n_0_0_171), .C2(n_0_0_139), .ZN(n_0_0_138));
   OAI21_X1 i_0_0_132 (.A(n_0_0_166), .B1(n_0_0), .B2(n_0_0_262), .ZN(n_0_0_139));
   INV_X1 i_0_0_133 (.A(n_0_0_140), .ZN(Sum[24]));
   AOI222_X1 i_0_0_134 (.A1(n_0_0_8), .A2(n_0_0_232), .B1(exp_Sum[1]), .B2(
      n_0_0_153), .C1(n_0_0_171), .C2(n_0_0_141), .ZN(n_0_0_140));
   XOR2_X1 i_0_0_135 (.A(n_0_0_166), .B(n_0_0_164), .Z(n_0_0_141));
   INV_X1 i_0_0_136 (.A(n_0_0_142), .ZN(Sum[25]));
   AOI222_X1 i_0_0_137 (.A1(n_0_0_9), .A2(n_0_0_232), .B1(exp_Sum[2]), .B2(
      n_0_0_153), .C1(n_0_0_171), .C2(n_0_0_143), .ZN(n_0_0_142));
   XOR2_X1 i_0_0_138 (.A(n_0_0_168), .B(n_0_0_163), .Z(n_0_0_143));
   INV_X1 i_0_0_139 (.A(n_0_0_144), .ZN(Sum[26]));
   AOI222_X1 i_0_0_140 (.A1(n_0_0_10), .A2(n_0_0_232), .B1(exp_Sum[3]), .B2(
      n_0_0_153), .C1(n_0_0_171), .C2(n_0_0_145), .ZN(n_0_0_144));
   XNOR2_X1 i_0_0_141 (.A(n_0_0_169), .B(n_0_0_162), .ZN(n_0_0_145));
   INV_X1 i_0_0_142 (.A(n_0_0_146), .ZN(Sum[27]));
   AOI222_X1 i_0_0_143 (.A1(n_0_0_11), .A2(n_0_0_232), .B1(exp_Sum[4]), .B2(
      n_0_0_153), .C1(n_0_0_171), .C2(n_0_0_147), .ZN(n_0_0_146));
   XOR2_X1 i_0_0_144 (.A(n_0_0_170), .B(n_0_0_161), .Z(n_0_0_147));
   OAI21_X1 i_0_0_145 (.A(n_0_0_148), .B1(n_0_0_267), .B2(n_0_0_154), .ZN(
      Sum[28]));
   AOI22_X1 i_0_0_146 (.A1(n_0_0_12), .A2(n_0_0_232), .B1(n_0_0_171), .B2(
      n_0_0_149), .ZN(n_0_0_148));
   OAI21_X1 i_0_0_147 (.A(n_0_0_159), .B1(n_0_0_267), .B2(n_0_0_160), .ZN(
      n_0_0_149));
   OAI211_X1 i_0_0_148 (.A(n_0_0_156), .B(n_0_0_150), .C1(n_0_0_268), .C2(
      n_0_0_151), .ZN(Sum[29]));
   NAND2_X1 i_0_0_149 (.A1(n_0_0_13), .A2(n_0_0_232), .ZN(n_0_0_150));
   AOI21_X1 i_0_0_150 (.A(n_0_0_153), .B1(n_0_0_171), .B2(n_0_0_159), .ZN(
      n_0_0_151));
   AOI22_X1 i_0_0_151 (.A1(n_0_0_156), .A2(n_0_0_155), .B1(exp_Sum[7]), .B2(
      n_0_0_152), .ZN(Sum[30]));
   AOI221_X1 i_0_0_152 (.A(n_0_0_153), .B1(n_0_0_171), .B2(n_0_0_157), .C1(
      n_0_0_563), .C2(n_0_0_232), .ZN(n_0_0_152));
   INV_X1 i_0_0_153 (.A(n_0_0_154), .ZN(n_0_0_153));
   NAND3_X1 i_0_0_154 (.A1(num_leading_zeros[4]), .A2(num_leading_zeros[3]), 
      .A3(n_0_0_230), .ZN(n_0_0_154));
   AOI21_X1 i_0_0_155 (.A(exp_Sum[7]), .B1(n_0_0_6), .B2(n_0_0_232), .ZN(
      n_0_0_155));
   NAND2_X1 i_0_0_156 (.A1(n_0_0_171), .A2(n_0_0_158), .ZN(n_0_0_156));
   INV_X1 i_0_0_157 (.A(n_0_0_158), .ZN(n_0_0_157));
   NOR2_X1 i_0_0_158 (.A1(exp_Sum[6]), .A2(n_0_0_159), .ZN(n_0_0_158));
   NAND2_X1 i_0_0_159 (.A1(n_0_0_267), .A2(n_0_0_160), .ZN(n_0_0_159));
   AOI22_X1 i_0_0_160 (.A1(n_0_0_129), .A2(exp_Sum[4]), .B1(n_0_0_170), .B2(
      n_0_0_161), .ZN(n_0_0_160));
   AOI22_X1 i_0_0_161 (.A1(n_0_3), .A2(n_0_0_265), .B1(n_0_0_169), .B2(n_0_0_162), 
      .ZN(n_0_0_161));
   OAI22_X1 i_0_0_162 (.A1(n_0_0_126), .A2(exp_Sum[2]), .B1(n_0_0_167), .B2(
      n_0_0_163), .ZN(n_0_0_162));
   AOI22_X1 i_0_0_163 (.A1(n_0_1), .A2(n_0_0_263), .B1(n_0_0_165), .B2(n_0_0_164), 
      .ZN(n_0_0_163));
   AOI22_X1 i_0_0_164 (.A1(n_0_1), .A2(n_0_0_263), .B1(n_0_0_125), .B2(
      exp_Sum[1]), .ZN(n_0_0_164));
   INV_X1 i_0_0_165 (.A(n_0_0_166), .ZN(n_0_0_165));
   NAND2_X1 i_0_0_166 (.A1(n_0_0), .A2(n_0_0_262), .ZN(n_0_0_166));
   INV_X1 i_0_0_167 (.A(n_0_0_168), .ZN(n_0_0_167));
   AOI22_X1 i_0_0_168 (.A1(n_0_2), .A2(n_0_0_264), .B1(n_0_0_126), .B2(
      exp_Sum[2]), .ZN(n_0_0_168));
   AOI22_X1 i_0_0_169 (.A1(n_0_3), .A2(n_0_0_265), .B1(n_0_0_128), .B2(
      exp_Sum[3]), .ZN(n_0_0_169));
   AOI22_X1 i_0_0_170 (.A1(n_0_0_129), .A2(exp_Sum[4]), .B1(n_0_4), .B2(
      n_0_0_266), .ZN(n_0_0_170));
   NOR2_X1 i_0_0_171 (.A1(n_0_5), .A2(n_0_0_228), .ZN(n_0_0_171));
   OAI21_X1 i_0_0_196 (.A(n_0_0_172), .B1(n_0_0_94), .B2(n_0_0_173), .ZN(Sum[31]));
   NAND2_X1 i_0_0_197 (.A1(A[31]), .A2(n_0_0_173), .ZN(n_0_0_172));
   AOI21_X1 i_0_0_198 (.A(n_0_0_396), .B1(n_48), .B2(n_0_0_174), .ZN(n_0_0_173));
   OAI22_X1 i_0_0_199 (.A1(n_0_0_613), .A2(A[22]), .B1(n_0_0_176), .B2(n_0_0_175), 
      .ZN(n_0_0_174));
   OAI22_X1 i_0_0_200 (.A1(B[21]), .A2(n_0_0_587), .B1(B[22]), .B2(n_0_0_588), 
      .ZN(n_0_0_175));
   AOI221_X1 i_0_0_201 (.A(n_0_0_177), .B1(B[21]), .B2(n_0_0_587), .C1(B[20]), 
      .C2(n_0_0_586), .ZN(n_0_0_176));
   AOI221_X1 i_0_0_202 (.A(n_0_0_178), .B1(n_0_0_611), .B2(A[19]), .C1(n_0_0_612), 
      .C2(A[20]), .ZN(n_0_0_177));
   AOI221_X1 i_0_0_203 (.A(n_0_0_179), .B1(B[19]), .B2(n_0_0_585), .C1(B[18]), 
      .C2(n_0_0_584), .ZN(n_0_0_178));
   AOI221_X1 i_0_0_204 (.A(n_0_0_180), .B1(n_0_0_609), .B2(A[17]), .C1(n_0_0_610), 
      .C2(A[18]), .ZN(n_0_0_179));
   AOI21_X1 i_0_0_205 (.A(n_0_0_181), .B1(B[17]), .B2(n_0_0_583), .ZN(n_0_0_180));
   AOI22_X1 i_0_0_206 (.A1(n_0_0_183), .A2(n_0_0_182), .B1(n_0_0_608), .B2(A[16]), 
      .ZN(n_0_0_181));
   AOI22_X1 i_0_0_207 (.A1(B[16]), .A2(n_0_0_582), .B1(B[15]), .B2(n_0_0_581), 
      .ZN(n_0_0_182));
   OAI221_X1 i_0_0_208 (.A(n_0_0_184), .B1(B[14]), .B2(n_0_0_580), .C1(B[15]), 
      .C2(n_0_0_581), .ZN(n_0_0_183));
   INV_X1 i_0_0_209 (.A(n_0_0_185), .ZN(n_0_0_184));
   AOI221_X1 i_0_0_210 (.A(n_0_0_186), .B1(B[13]), .B2(n_0_0_579), .C1(B[14]), 
      .C2(n_0_0_580), .ZN(n_0_0_185));
   AOI21_X1 i_0_0_211 (.A(n_0_0_187), .B1(n_0_0_607), .B2(A[13]), .ZN(n_0_0_186));
   AOI22_X1 i_0_0_212 (.A1(n_0_0_189), .A2(n_0_0_188), .B1(B[12]), .B2(n_0_0_578), 
      .ZN(n_0_0_187));
   AOI22_X1 i_0_0_213 (.A1(n_0_0_606), .A2(A[12]), .B1(n_0_0_605), .B2(A[11]), 
      .ZN(n_0_0_188));
   OAI221_X1 i_0_0_214 (.A(n_0_0_190), .B1(n_0_0_604), .B2(A[10]), .C1(n_0_0_605), 
      .C2(A[11]), .ZN(n_0_0_189));
   INV_X1 i_0_0_215 (.A(n_0_0_191), .ZN(n_0_0_190));
   AOI221_X1 i_0_0_216 (.A(n_0_0_362), .B1(n_0_0_603), .B2(A[9]), .C1(n_0_0_604), 
      .C2(A[10]), .ZN(n_0_0_191));
   AOI21_X1 i_0_0_172 (.A(n_0_0_203), .B1(n_0_0_274), .B2(n_0_0_231), .ZN(
      mant_A[1]));
   NOR2_X1 i_0_0_173 (.A1(n_0_6), .A2(n_0_0_231), .ZN(n_0_0_203));
   AOI21_X1 i_0_0_174 (.A(n_0_0_204), .B1(n_0_0_279), .B2(n_0_0_231), .ZN(
      mant_A[2]));
   NOR2_X1 i_0_0_175 (.A1(n_0_7), .A2(n_0_0_231), .ZN(n_0_0_204));
   AOI21_X1 i_0_0_176 (.A(n_0_0_205), .B1(n_0_0_284), .B2(n_0_0_231), .ZN(
      mant_A[3]));
   NOR2_X1 i_0_0_177 (.A1(n_0_8), .A2(n_0_0_231), .ZN(n_0_0_205));
   AOI21_X1 i_0_0_178 (.A(n_0_0_206), .B1(n_0_0_290), .B2(n_0_0_231), .ZN(
      mant_A[4]));
   NOR2_X1 i_0_0_179 (.A1(n_0_9), .A2(n_0_0_231), .ZN(n_0_0_206));
   AOI21_X1 i_0_0_180 (.A(n_0_0_207), .B1(n_0_0_295), .B2(n_0_0_231), .ZN(
      mant_A[5]));
   NOR2_X1 i_0_0_181 (.A1(n_0_10), .A2(n_0_0_231), .ZN(n_0_0_207));
   AOI21_X1 i_0_0_182 (.A(n_0_0_208), .B1(n_0_0_300), .B2(n_0_0_231), .ZN(
      mant_A[6]));
   NOR2_X1 i_0_0_183 (.A1(n_0_11), .A2(n_0_0_231), .ZN(n_0_0_208));
   AOI21_X1 i_0_0_184 (.A(n_0_0_209), .B1(n_0_0_366), .B2(n_0_0_231), .ZN(
      mant_A[7]));
   NOR2_X1 i_0_0_185 (.A1(n_0_12), .A2(n_0_0_231), .ZN(n_0_0_209));
   AOI21_X1 i_0_0_186 (.A(n_0_0_210), .B1(n_0_0_311), .B2(n_0_0_231), .ZN(
      mant_A[8]));
   NOR2_X1 i_0_0_187 (.A1(n_0_13), .A2(n_0_0_231), .ZN(n_0_0_210));
   AOI21_X1 i_0_0_188 (.A(n_0_0_211), .B1(n_0_0_317), .B2(n_0_0_231), .ZN(
      mant_A[9]));
   NOR2_X1 i_0_0_189 (.A1(n_0_14), .A2(n_0_0_231), .ZN(n_0_0_211));
   AOI21_X1 i_0_0_190 (.A(n_0_0_212), .B1(n_0_0_320), .B2(n_0_0_231), .ZN(
      mant_A[10]));
   NOR2_X1 i_0_0_191 (.A1(n_0_15), .A2(n_0_0_231), .ZN(n_0_0_212));
   AOI21_X1 i_0_0_192 (.A(n_0_0_213), .B1(n_0_0_328), .B2(n_0_0_231), .ZN(
      mant_A[11]));
   NOR2_X1 i_0_0_193 (.A1(n_0_16), .A2(n_0_0_231), .ZN(n_0_0_213));
   AOI21_X1 i_0_0_194 (.A(n_0_0_214), .B1(n_0_0_334), .B2(n_0_0_231), .ZN(
      mant_A[12]));
   NOR2_X1 i_0_0_195 (.A1(n_0_17), .A2(n_0_0_231), .ZN(n_0_0_214));
   AOI21_X1 i_0_0_217 (.A(n_0_0_215), .B1(n_0_0_337), .B2(n_0_0_231), .ZN(
      mant_A[13]));
   NOR2_X1 i_0_0_218 (.A1(n_0_18), .A2(n_0_0_231), .ZN(n_0_0_215));
   AOI21_X1 i_0_0_219 (.A(n_0_0_216), .B1(n_0_0_342), .B2(n_0_0_231), .ZN(
      mant_A[14]));
   NOR2_X1 i_0_0_220 (.A1(n_0_19), .A2(n_0_0_231), .ZN(n_0_0_216));
   AOI21_X1 i_0_0_221 (.A(n_0_0_217), .B1(n_0_0_346), .B2(n_0_0_231), .ZN(
      mant_A[15]));
   NOR2_X1 i_0_0_222 (.A1(n_0_20), .A2(n_0_0_231), .ZN(n_0_0_217));
   AOI21_X1 i_0_0_223 (.A(n_0_0_218), .B1(n_0_0_356), .B2(n_0_0_231), .ZN(
      mant_A[16]));
   NOR2_X1 i_0_0_224 (.A1(n_0_21), .A2(n_0_0_231), .ZN(n_0_0_218));
   AOI21_X1 i_0_0_225 (.A(n_0_0_219), .B1(n_0_0_359), .B2(n_0_0_231), .ZN(
      mant_A[17]));
   NOR2_X1 i_0_0_226 (.A1(n_0_22), .A2(n_0_0_231), .ZN(n_0_0_219));
   AOI21_X1 i_0_0_227 (.A(n_0_0_220), .B1(n_0_0_363), .B2(n_0_0_231), .ZN(
      mant_A[18]));
   NOR2_X1 i_0_0_228 (.A1(n_0_23), .A2(n_0_0_231), .ZN(n_0_0_220));
   AOI21_X1 i_0_0_229 (.A(n_0_0_221), .B1(n_0_0_367), .B2(n_0_0_231), .ZN(
      mant_A[19]));
   NOR2_X1 i_0_0_230 (.A1(n_0_24), .A2(n_0_0_231), .ZN(n_0_0_221));
   AOI21_X1 i_0_0_231 (.A(n_0_0_222), .B1(n_0_0_376), .B2(n_0_0_231), .ZN(
      mant_A[20]));
   NOR2_X1 i_0_0_232 (.A1(n_0_25), .A2(n_0_0_231), .ZN(n_0_0_222));
   AOI21_X1 i_0_0_233 (.A(n_0_0_223), .B1(n_0_0_379), .B2(n_0_0_231), .ZN(
      mant_A[21]));
   NOR2_X1 i_0_0_234 (.A1(n_0_26), .A2(n_0_0_231), .ZN(n_0_0_223));
   AOI21_X1 i_0_0_235 (.A(n_0_0_224), .B1(n_0_0_381), .B2(n_0_0_231), .ZN(
      mant_A[22]));
   NOR2_X1 i_0_0_236 (.A1(n_0_27), .A2(n_0_0_231), .ZN(n_0_0_224));
   AOI22_X1 i_0_0_237 (.A1(n_0_0_564), .A2(n_0_0_230), .B1(n_0_0_396), .B2(
      n_0_0_232), .ZN(mant_A[23]));
   AND2_X1 i_0_0_238 (.A1(n_0_29), .A2(n_0_0_230), .ZN(mant_A[31]));
   NOR2_X1 i_0_0_239 (.A1(n_0_0_233), .A2(n_0_0_225), .ZN(overflow));
   NAND4_X1 i_0_0_240 (.A1(n_24), .A2(exp_Sum[7]), .A3(exp_Sum[6]), .A4(
      n_0_0_226), .ZN(n_0_0_225));
   NOR4_X1 i_0_0_241 (.A1(exp_Sum[0]), .A2(n_0_0_227), .A3(n_0_0_267), .A4(
      n_0_0_266), .ZN(n_0_0_226));
   NAND3_X1 i_0_0_242 (.A1(exp_Sum[3]), .A2(exp_Sum[2]), .A3(exp_Sum[1]), 
      .ZN(n_0_0_227));
   AND2_X1 i_0_0_278 (.A1(n_0_5), .A2(n_0_0_229), .ZN(underflow));
   INV_X1 i_0_0_243 (.A(n_0_0_229), .ZN(n_0_0_228));
   AOI21_X1 i_0_0_244 (.A(n_0_0_231), .B1(num_leading_zeros[4]), .B2(
      num_leading_zeros[3]), .ZN(n_0_0_229));
   INV_X1 i_0_0_245 (.A(n_0_0_231), .ZN(n_0_0_230));
   OAI21_X1 i_0_0_246 (.A(n_0_0_233), .B1(n_0_0_246), .B2(n_0_0_234), .ZN(
      n_0_0_231));
   INV_X1 i_0_0_247 (.A(n_0_0_233), .ZN(n_0_0_232));
   XNOR2_X1 i_0_0_248 (.A(n_0_0_94), .B(A[31]), .ZN(n_0_0_233));
   NAND4_X1 i_0_0_249 (.A1(n_0_0_253), .A2(n_0_0_235), .A3(n_0_0_236), .A4(
      n_0_0_238), .ZN(n_0_0_234));
   AOI221_X1 i_0_0_250 (.A(n_0_0_259), .B1(n_33), .B2(n_0_0_317), .C1(n_28), 
      .C2(n_0_0_284), .ZN(n_0_0_235));
   AOI221_X1 i_0_0_251 (.A(n_0_0_237), .B1(n_0_0_458), .B2(n_0_42), .C1(n_37), 
      .C2(n_0_0_337), .ZN(n_0_0_236));
   OAI222_X1 i_0_0_252 (.A1(n_28), .A2(n_0_0_284), .B1(n_0_0_406), .B2(n_0_31), 
      .C1(n_0_0_416), .C2(n_0_33), .ZN(n_0_0_237));
   NOR4_X1 i_0_0_253 (.A1(n_0_0_260), .A2(n_0_0_245), .A3(n_0_0_244), .A4(
      n_0_0_239), .ZN(n_0_0_238));
   NAND4_X1 i_0_0_254 (.A1(n_0_0_243), .A2(n_0_0_242), .A3(n_0_0_241), .A4(
      n_0_0_240), .ZN(n_0_0_239));
   AOI22_X1 i_0_0_255 (.A1(n_0_0_467), .A2(n_0_44), .B1(n_0_0_461), .B2(n_0_43), 
      .ZN(n_0_0_240));
   AOI221_X1 i_0_0_256 (.A(n_0_0_255), .B1(n_0_0_477), .B2(n_0_46), .C1(
      n_0_0_473), .C2(n_0_45), .ZN(n_0_0_241));
   AOI22_X1 i_0_0_257 (.A1(n_39), .A2(n_0_0_346), .B1(n_38), .B2(n_0_0_342), 
      .ZN(n_0_0_242));
   AOI22_X1 i_0_0_258 (.A1(n_42), .A2(n_0_0_363), .B1(n_0_0_481), .B2(n_0_47), 
      .ZN(n_0_0_243));
   OAI21_X1 i_0_0_259 (.A(n_0_0_261), .B1(n_29), .B2(n_0_0_290), .ZN(n_0_0_244));
   OAI221_X1 i_0_0_260 (.A(n_0_0_254), .B1(n_27), .B2(n_0_0_279), .C1(n_26), 
      .C2(n_0_0_274), .ZN(n_0_0_245));
   OAI221_X1 i_0_0_261 (.A(n_0_0_247), .B1(n_0_0_397), .B2(mant_A[0]), .C1(n_25), 
      .C2(n_0_0_269), .ZN(n_0_0_246));
   AOI221_X1 i_0_0_262 (.A(n_0_0_248), .B1(n_0_0_550), .B2(n_0_34), .C1(n_47), 
      .C2(n_0_0_295), .ZN(n_0_0_247));
   OAI211_X1 i_0_0_263 (.A(n_0_0_252), .B(n_0_0_249), .C1(n_0_0_437), .C2(n_0_37), 
      .ZN(n_0_0_248));
   AOI221_X1 i_0_0_264 (.A(n_0_0_250), .B1(n_34), .B2(n_0_0_320), .C1(n_0_0_437), 
      .C2(n_0_37), .ZN(n_0_0_249));
   OAI221_X1 i_0_0_265 (.A(n_0_0_251), .B1(n_0_0_487), .B2(n_0_48), .C1(n_43), 
      .C2(n_0_0_367), .ZN(n_0_0_250));
   AOI222_X1 i_0_0_266 (.A1(n_41), .A2(n_0_0_359), .B1(n_40), .B2(n_0_0_356), 
      .C1(n_0_0_426), .C2(n_0_35), .ZN(n_0_0_251));
   AOI22_X1 i_0_0_267 (.A1(n_30), .A2(n_0_0_300), .B1(n_0_0_446), .B2(n_0_39), 
      .ZN(n_0_0_252));
   OAI22_X1 i_0_0_268 (.A1(n_0_0_431), .A2(n_0_0_366), .B1(n_31), .B2(n_0_36), 
      .ZN(n_0_0_253));
   AOI22_X1 i_0_0_269 (.A1(n_0_0_451), .A2(n_0_40), .B1(n_35), .B2(n_0_0_328), 
      .ZN(n_0_0_254));
   NAND3_X1 i_0_0_270 (.A1(n_0_0_257), .A2(n_0_0_256), .A3(n_0_0_258), .ZN(
      n_0_0_255));
   AOI211_X1 i_0_0_271 (.A(n_0_0_506), .B(n_0_0_517), .C1(n_44), .C2(n_0_0_376), 
      .ZN(n_0_0_256));
   XOR2_X1 i_0_0_272 (.A(n_46), .B(n_0_0_381), .Z(n_0_0_257));
   AOI222_X1 i_0_0_273 (.A1(n_0_0_501), .A2(n_0_50), .B1(n_0_0_496), .B2(n_0_49), 
      .C1(n_45), .C2(n_0_0_379), .ZN(n_0_0_258));
   NOR2_X1 i_0_0_274 (.A1(n_33), .A2(n_0_0_317), .ZN(n_0_0_259));
   XOR2_X1 i_0_0_275 (.A(n_36), .B(n_0_41), .Z(n_0_0_260));
   NAND2_X1 i_0_0_276 (.A1(n_26), .A2(n_0_0_274), .ZN(n_0_0_261));
   INV_X1 i_0_0_277 (.A(n_0_0_262), .ZN(exp_Sum[0]));
   AOI22_X1 i_0_0_279 (.A1(B[23]), .A2(n_0_0_396), .B1(A[23]), .B2(n_0_52), 
      .ZN(n_0_0_262));
   INV_X1 i_0_0_280 (.A(n_0_0_263), .ZN(exp_Sum[1]));
   AOI22_X1 i_0_0_281 (.A1(B[24]), .A2(n_0_0_396), .B1(A[24]), .B2(n_0_52), 
      .ZN(n_0_0_263));
   INV_X1 i_0_0_282 (.A(n_0_0_264), .ZN(exp_Sum[2]));
   AOI22_X1 i_0_0_283 (.A1(B[25]), .A2(n_0_0_396), .B1(A[25]), .B2(n_0_52), 
      .ZN(n_0_0_264));
   INV_X1 i_0_0_284 (.A(n_0_0_265), .ZN(exp_Sum[3]));
   AOI22_X1 i_0_0_285 (.A1(B[26]), .A2(n_0_0_396), .B1(A[26]), .B2(n_0_52), 
      .ZN(n_0_0_265));
   INV_X1 i_0_0_286 (.A(n_0_0_266), .ZN(exp_Sum[4]));
   AOI22_X1 i_0_0_287 (.A1(B[27]), .A2(n_0_0_396), .B1(A[27]), .B2(n_0_52), 
      .ZN(n_0_0_266));
   INV_X1 i_0_0_288 (.A(n_0_0_267), .ZN(exp_Sum[5]));
   AOI22_X1 i_0_0_289 (.A1(B[28]), .A2(n_0_0_396), .B1(A[28]), .B2(n_0_52), 
      .ZN(n_0_0_267));
   INV_X1 i_0_0_290 (.A(n_0_0_268), .ZN(exp_Sum[6]));
   AOI22_X1 i_0_0_291 (.A1(B[29]), .A2(n_0_0_396), .B1(A[29]), .B2(n_0_52), 
      .ZN(n_0_0_268));
   INV_X1 i_0_0_292 (.A(n_0_0_269), .ZN(mant_A[0]));
   AOI221_X1 i_0_0_293 (.A(n_0_0_270), .B1(A[0]), .B2(n_0_52), .C1(n_0_0_390), 
      .C2(n_0_0_275), .ZN(n_0_0_269));
   AOI221_X1 i_0_0_294 (.A(n_0_0_471), .B1(n_0_0_470), .B2(n_0_0_271), .C1(
      n_0_0_450), .C2(n_0_0_281), .ZN(n_0_0_270));
   AOI221_X1 i_0_0_295 (.A(n_0_0_272), .B1(A[8]), .B2(n_0_0_388), .C1(A[16]), 
      .C2(n_0_0_289), .ZN(n_0_0_271));
   INV_X1 i_0_0_296 (.A(n_0_0_273), .ZN(n_0_0_272));
   AOI22_X1 i_0_0_297 (.A1(n_0_0_441), .A2(n_0_0_293), .B1(A[0]), .B2(n_0_0_422), 
      .ZN(n_0_0_273));
   INV_X1 i_0_0_333 (.A(n_0_0_274), .ZN(n_0_30));
   AOI222_X1 i_0_0_298 (.A1(n_0_0_390), .A2(n_0_0_280), .B1(A[1]), .B2(n_0_52), 
      .C1(n_0_0_484), .C2(n_0_0_275), .ZN(n_0_0_274));
   AOI22_X1 i_0_0_299 (.A1(n_0_0_450), .A2(n_0_0_286), .B1(n_0_0_470), .B2(
      n_0_0_276), .ZN(n_0_0_275));
   AOI221_X1 i_0_0_300 (.A(n_0_0_277), .B1(A[17]), .B2(n_0_0_289), .C1(n_0_0_441), 
      .C2(n_0_0_298), .ZN(n_0_0_276));
   OAI21_X1 i_0_0_301 (.A(n_0_0_278), .B1(n_0_0_198), .B2(n_0_0_421), .ZN(
      n_0_0_277));
   NAND2_X1 i_0_0_302 (.A1(A[9]), .A2(n_0_0_388), .ZN(n_0_0_278));
   INV_X1 i_0_0_303 (.A(n_0_0_279), .ZN(n_0_31));
   AOI222_X1 i_0_0_304 (.A1(n_0_0_484), .A2(n_0_0_280), .B1(A[2]), .B2(n_0_52), 
      .C1(n_0_0_390), .C2(n_0_0_285), .ZN(n_0_0_279));
   AOI22_X1 i_0_0_305 (.A1(n_0_0_470), .A2(n_0_0_281), .B1(n_0_0_450), .B2(
      n_0_0_292), .ZN(n_0_0_280));
   AOI221_X1 i_0_0_306 (.A(n_0_0_282), .B1(A[18]), .B2(n_0_0_289), .C1(A[2]), 
      .C2(n_0_0_422), .ZN(n_0_0_281));
   INV_X1 i_0_0_307 (.A(n_0_0_283), .ZN(n_0_0_282));
   AOI22_X1 i_0_0_308 (.A1(n_0_0_441), .A2(n_0_0_303), .B1(A[10]), .B2(n_0_0_388), 
      .ZN(n_0_0_283));
   INV_X1 i_0_0_345 (.A(n_0_0_284), .ZN(n_0_32));
   AOI222_X1 i_0_0_309 (.A1(n_0_0_390), .A2(n_0_0_291), .B1(A[3]), .B2(n_0_52), 
      .C1(n_0_0_484), .C2(n_0_0_285), .ZN(n_0_0_284));
   AOI22_X1 i_0_0_310 (.A1(n_0_0_470), .A2(n_0_0_286), .B1(n_0_0_450), .B2(
      n_0_0_297), .ZN(n_0_0_285));
   AOI221_X1 i_0_0_311 (.A(n_0_0_287), .B1(A[19]), .B2(n_0_0_289), .C1(A[3]), 
      .C2(n_0_0_422), .ZN(n_0_0_286));
   INV_X1 i_0_0_312 (.A(n_0_0_288), .ZN(n_0_0_287));
   AOI22_X1 i_0_0_313 (.A1(n_0_0_441), .A2(n_0_0_424), .B1(A[11]), .B2(n_0_0_388), 
      .ZN(n_0_0_288));
   NOR3_X1 i_0_0_314 (.A1(n_0_0_439), .A2(n_0_0_435), .A3(n_0_0_441), .ZN(
      n_0_0_289));
   INV_X1 i_0_0_315 (.A(n_0_0_290), .ZN(n_0_33));
   AOI222_X1 i_0_0_316 (.A1(n_0_0_390), .A2(n_0_0_296), .B1(A[4]), .B2(n_0_52), 
      .C1(n_0_0_484), .C2(n_0_0_291), .ZN(n_0_0_290));
   AOI22_X1 i_0_0_317 (.A1(n_0_0_470), .A2(n_0_0_292), .B1(n_0_0_450), .B2(
      n_0_0_302), .ZN(n_0_0_291));
   AOI222_X1 i_0_0_318 (.A1(A[16]), .A2(n_0_0_389), .B1(A[8]), .B2(n_0_0_394), 
      .C1(n_0_0_442), .C2(n_0_0_293), .ZN(n_0_0_292));
   OAI21_X1 i_0_0_319 (.A(n_0_0_294), .B1(n_0_0_306), .B2(n_0_0_430), .ZN(
      n_0_0_293));
   AOI22_X1 i_0_0_320 (.A1(A[12]), .A2(n_0_0_433), .B1(A[20]), .B2(n_0_0_305), 
      .ZN(n_0_0_294));
   INV_X1 i_0_0_321 (.A(n_0_0_295), .ZN(n_0_34));
   AOI222_X1 i_0_0_322 (.A1(n_0_0_390), .A2(n_0_0_301), .B1(A[5]), .B2(n_0_52), 
      .C1(n_0_0_484), .C2(n_0_0_296), .ZN(n_0_0_295));
   AOI22_X1 i_0_0_323 (.A1(n_0_0_470), .A2(n_0_0_297), .B1(n_0_0_450), .B2(
      n_0_0_423), .ZN(n_0_0_296));
   AOI222_X1 i_0_0_324 (.A1(A[17]), .A2(n_0_0_389), .B1(A[9]), .B2(n_0_0_394), 
      .C1(n_0_0_442), .C2(n_0_0_298), .ZN(n_0_0_297));
   OAI21_X1 i_0_0_325 (.A(n_0_0_299), .B1(n_0_0_307), .B2(n_0_0_430), .ZN(
      n_0_0_298));
   AOI22_X1 i_0_0_326 (.A1(A[13]), .A2(n_0_0_433), .B1(A[21]), .B2(n_0_0_305), 
      .ZN(n_0_0_299));
   INV_X1 i_0_0_327 (.A(n_0_0_300), .ZN(n_0_35));
   AOI222_X1 i_0_0_328 (.A1(A[6]), .A2(n_0_52), .B1(n_0_0_390), .B2(n_0_0_391), 
      .C1(n_0_0_484), .C2(n_0_0_301), .ZN(n_0_0_300));
   AOI22_X1 i_0_0_329 (.A1(n_0_0_470), .A2(n_0_0_302), .B1(n_0_0_450), .B2(
      n_0_0_374), .ZN(n_0_0_301));
   AOI222_X1 i_0_0_330 (.A1(A[18]), .A2(n_0_0_389), .B1(A[10]), .B2(n_0_0_394), 
      .C1(n_0_0_442), .C2(n_0_0_303), .ZN(n_0_0_302));
   OAI21_X1 i_0_0_331 (.A(n_0_0_304), .B1(n_0_0_309), .B2(n_0_0_430), .ZN(
      n_0_0_303));
   AOI22_X1 i_0_0_332 (.A1(A[14]), .A2(n_0_0_433), .B1(A[22]), .B2(n_0_0_305), 
      .ZN(n_0_0_304));
   NOR2_X1 i_0_0_334 (.A1(n_0_0_439), .A2(n_0_0_435), .ZN(n_0_0_305));
   INV_X1 i_0_0_335 (.A(n_0_0_311), .ZN(n_0_37));
   AOI222_X1 i_0_0_336 (.A1(n_0_0_390), .A2(n_0_0_318), .B1(A[8]), .B2(n_0_52), 
      .C1(n_0_0_484), .C2(n_0_0_369), .ZN(n_0_0_311));
   INV_X1 i_0_0_337 (.A(n_0_0_317), .ZN(n_0_38));
   AOI222_X1 i_0_0_338 (.A1(n_0_0_390), .A2(n_0_0_321), .B1(A[9]), .B2(n_0_52), 
      .C1(n_0_0_484), .C2(n_0_0_318), .ZN(n_0_0_317));
   AOI22_X1 i_0_0_339 (.A1(n_0_0_470), .A2(n_0_0_392), .B1(n_0_0_450), .B2(
      n_0_0_331), .ZN(n_0_0_318));
   INV_X1 i_0_0_340 (.A(n_0_0_320), .ZN(n_0_39));
   AOI222_X1 i_0_0_341 (.A1(n_0_0_390), .A2(n_0_0_329), .B1(A[10]), .B2(n_0_52), 
      .C1(n_0_0_484), .C2(n_0_0_321), .ZN(n_0_0_320));
   AOI21_X1 i_0_0_342 (.A(n_0_0_322), .B1(n_0_0_450), .B2(n_0_0_336), .ZN(
      n_0_0_321));
   NOR2_X1 i_0_0_343 (.A1(n_0_0_450), .A2(n_0_0_384), .ZN(n_0_0_322));
   INV_X1 i_0_0_344 (.A(n_0_0_328), .ZN(n_0_40));
   AOI222_X1 i_0_0_346 (.A1(n_0_0_484), .A2(n_0_0_329), .B1(A[11]), .B2(n_0_52), 
      .C1(n_0_0_390), .C2(n_0_0_335), .ZN(n_0_0_328));
   OAI21_X1 i_0_0_347 (.A(n_0_0_330), .B1(n_0_0_450), .B2(n_0_0_331), .ZN(
      n_0_0_329));
   NAND2_X1 i_0_0_348 (.A1(n_0_0_450), .A2(n_0_0_340), .ZN(n_0_0_330));
   INV_X1 i_0_0_349 (.A(n_0_0_332), .ZN(n_0_0_331));
   AOI22_X1 i_0_0_350 (.A1(n_0_0_442), .A2(n_0_0_428), .B1(n_0_0_441), .B2(
      n_0_0_351), .ZN(n_0_0_332));
   INV_X1 i_0_0_351 (.A(n_0_0_334), .ZN(n_0_41));
   AOI222_X1 i_0_0_352 (.A1(n_0_0_390), .A2(n_0_0_338), .B1(A[12]), .B2(n_0_52), 
      .C1(n_0_0_484), .C2(n_0_0_335), .ZN(n_0_0_334));
   AOI22_X1 i_0_0_353 (.A1(n_0_0_470), .A2(n_0_0_336), .B1(n_0_0_450), .B2(
      n_0_0_344), .ZN(n_0_0_335));
   AOI222_X1 i_0_0_354 (.A1(A[16]), .A2(n_0_0_394), .B1(A[12]), .B2(n_0_0_422), 
      .C1(A[20]), .C2(n_0_0_388), .ZN(n_0_0_336));
   INV_X1 i_0_0_355 (.A(n_0_0_337), .ZN(n_0_42));
   AOI222_X1 i_0_0_356 (.A1(n_0_0_390), .A2(n_0_0_343), .B1(A[13]), .B2(n_0_52), 
      .C1(n_0_0_484), .C2(n_0_0_338), .ZN(n_0_0_337));
   INV_X1 i_0_0_357 (.A(n_0_0_339), .ZN(n_0_0_338));
   AOI22_X1 i_0_0_358 (.A1(n_0_0_450), .A2(n_0_0_350), .B1(n_0_0_470), .B2(
      n_0_0_340), .ZN(n_0_0_339));
   OAI21_X1 i_0_0_359 (.A(n_0_0_341), .B1(n_0_0_579), .B2(n_0_0_421), .ZN(
      n_0_0_340));
   AOI22_X1 i_0_0_360 (.A1(A[21]), .A2(n_0_0_388), .B1(A[17]), .B2(n_0_0_394), 
      .ZN(n_0_0_341));
   INV_X1 i_0_0_361 (.A(n_0_0_342), .ZN(n_0_43));
   AOI222_X1 i_0_0_362 (.A1(A[14]), .A2(n_0_52), .B1(n_0_0_390), .B2(n_0_0_347), 
      .C1(n_0_0_484), .C2(n_0_0_343), .ZN(n_0_0_342));
   AOI22_X1 i_0_0_363 (.A1(n_0_0_450), .A2(n_0_0_358), .B1(n_0_0_470), .B2(
      n_0_0_344), .ZN(n_0_0_343));
   AOI222_X1 i_0_0_364 (.A1(A[22]), .A2(n_0_0_388), .B1(A[14]), .B2(n_0_0_422), 
      .C1(A[18]), .C2(n_0_0_394), .ZN(n_0_0_344));
   INV_X1 i_0_0_365 (.A(n_0_0_346), .ZN(n_0_44));
   AOI222_X1 i_0_0_366 (.A1(n_0_0_484), .A2(n_0_0_347), .B1(A[15]), .B2(n_0_52), 
      .C1(n_0_0_390), .C2(n_0_0_357), .ZN(n_0_0_346));
   INV_X1 i_0_0_367 (.A(n_0_0_348), .ZN(n_0_0_347));
   AOI21_X1 i_0_0_368 (.A(n_0_0_349), .B1(n_0_0_470), .B2(n_0_0_350), .ZN(
      n_0_0_348));
   NOR3_X1 i_0_0_369 (.A1(n_0_0_430), .A2(n_0_0_395), .A3(n_0_0_470), .ZN(
      n_0_0_349));
   OAI21_X1 i_0_0_370 (.A(n_0_0_355), .B1(n_0_0_441), .B2(n_0_0_351), .ZN(
      n_0_0_350));
   AND2_X1 i_0_0_371 (.A1(n_0_0_434), .A2(n_0_0_425), .ZN(n_0_0_351));
   NAND2_X1 i_0_0_372 (.A1(A[19]), .A2(n_0_0_394), .ZN(n_0_0_355));
   INV_X1 i_0_0_373 (.A(n_0_0_356), .ZN(n_0_45));
   AOI222_X1 i_0_0_374 (.A1(n_0_0_390), .A2(n_0_0_360), .B1(A[16]), .B2(n_0_52), 
      .C1(n_0_0_484), .C2(n_0_0_357), .ZN(n_0_0_356));
   AOI22_X1 i_0_0_375 (.A1(n_0_0_450), .A2(n_0_0_365), .B1(n_0_0_470), .B2(
      n_0_0_358), .ZN(n_0_0_357));
   AOI22_X1 i_0_0_376 (.A1(A[16]), .A2(n_0_0_422), .B1(A[20]), .B2(n_0_0_394), 
      .ZN(n_0_0_358));
   INV_X1 i_0_0_377 (.A(n_0_0_359), .ZN(n_0_46));
   AOI222_X1 i_0_0_378 (.A1(n_0_0_484), .A2(n_0_0_360), .B1(A[17]), .B2(n_0_52), 
      .C1(n_0_0_390), .C2(n_0_0_364), .ZN(n_0_0_359));
   AOI221_X1 i_0_0_379 (.A(n_0_0_430), .B1(n_0_0_470), .B2(n_0_0_395), .C1(
      n_0_0_450), .C2(n_0_0_372), .ZN(n_0_0_360));
   INV_X1 i_0_0_380 (.A(n_0_0_363), .ZN(n_0_47));
   AOI222_X1 i_0_0_381 (.A1(A[18]), .A2(n_0_52), .B1(n_0_0_371), .B2(n_0_0_390), 
      .C1(n_0_0_484), .C2(n_0_0_364), .ZN(n_0_0_363));
   OAI22_X1 i_0_0_382 (.A1(n_0_0_586), .A2(n_0_0_373), .B1(n_0_0_450), .B2(
      n_0_0_365), .ZN(n_0_0_364));
   AOI22_X1 i_0_0_383 (.A1(A[18]), .A2(n_0_0_422), .B1(A[22]), .B2(n_0_0_394), 
      .ZN(n_0_0_365));
   INV_X1 i_0_0_384 (.A(n_0_0_367), .ZN(n_0_48));
   AOI221_X1 i_0_0_385 (.A(n_0_0_368), .B1(n_0_0_484), .B2(n_0_0_371), .C1(A[19]), 
      .C2(n_0_52), .ZN(n_0_0_367));
   AND3_X1 i_0_0_386 (.A1(n_0_0_422), .A2(n_0_0_370), .A3(n_0_0_390), .ZN(
      n_0_0_368));
   OAI22_X1 i_0_0_387 (.A1(n_0_0_588), .A2(n_0_0_470), .B1(n_0_0_586), .B2(
      n_0_0_450), .ZN(n_0_0_370));
   OAI33_X1 i_0_0_388 (.A1(n_0_0_470), .A2(n_0_0_421), .A3(n_0_0_587), .B1(
      n_0_0_430), .B2(n_0_0_372), .B3(n_0_0_450), .ZN(n_0_0_371));
   NOR2_X1 i_0_0_389 (.A1(A[19]), .A2(n_0_0_441), .ZN(n_0_0_372));
   NAND2_X1 i_0_0_390 (.A1(n_0_0_450), .A2(n_0_0_422), .ZN(n_0_0_373));
   INV_X1 i_0_0_391 (.A(n_0_0_376), .ZN(n_0_49));
   AOI22_X1 i_0_0_392 (.A1(A[20]), .A2(n_0_52), .B1(n_0_0_382), .B2(n_0_0_377), 
      .ZN(n_0_0_376));
   AOI21_X1 i_0_0_393 (.A(n_0_0_378), .B1(n_0_0_587), .B2(n_0_0_470), .ZN(
      n_0_0_377));
   AOI21_X1 i_0_0_394 (.A(n_0_0_539), .B1(A[22]), .B2(n_0_0_450), .ZN(n_0_0_378));
   INV_X1 i_0_0_395 (.A(n_0_0_379), .ZN(n_0_50));
   AOI22_X1 i_0_0_396 (.A1(A[21]), .A2(n_0_52), .B1(n_0_0_382), .B2(n_0_0_380), 
      .ZN(n_0_0_379));
   AOI21_X1 i_0_0_397 (.A(n_0_0_597), .B1(n_0_0_588), .B2(n_0_0_599), .ZN(
      n_0_0_380));
   INV_X1 i_0_0_461 (.A(n_0_0_381), .ZN(n_0_51));
   AOI22_X1 i_0_0_398 (.A1(A[22]), .A2(n_0_52), .B1(n_0_0_470), .B2(n_0_0_382), 
      .ZN(n_0_0_381));
   AND2_X1 i_0_0_399 (.A1(n_0_0_422), .A2(n_0_0_492), .ZN(n_0_0_382));
   INV_X1 i_0_0_400 (.A(n_0_52), .ZN(n_0_0_396));
   INV_X1 i_0_0_401 (.A(n_0_0_397), .ZN(n_25));
   AOI221_X1 i_0_0_402 (.A(n_0_0_398), .B1(B[0]), .B2(n_48), .C1(n_0_0_600), 
      .C2(n_0_0_402), .ZN(n_0_0_397));
   AOI221_X1 i_0_0_403 (.A(n_0_0_559), .B1(n_0_0_400), .B2(n_0_0_399), .C1(
      n_0_0_510), .C2(n_0_0_408), .ZN(n_0_0_398));
   AOI222_X1 i_0_0_404 (.A1(B[8]), .A2(n_0_0_572), .B1(B[0]), .B2(n_0_0_515), 
      .C1(n_0_0_594), .C2(n_0_0_419), .ZN(n_0_0_399));
   AOI21_X1 i_0_0_405 (.A(n_0_0_598), .B1(B[16]), .B2(n_0_0_414), .ZN(n_0_0_400));
   OAI21_X1 i_0_0_406 (.A(n_0_0_401), .B1(n_0_0_200), .B2(n_0_0_617), .ZN(n_26));
   AOI22_X1 i_0_0_407 (.A1(n_0_0_558), .A2(n_0_0_402), .B1(n_0_0_600), .B2(
      n_0_0_407), .ZN(n_0_0_401));
   AOI22_X1 i_0_0_408 (.A1(n_0_0_598), .A2(n_0_0_412), .B1(n_0_0_597), .B2(
      n_0_0_403), .ZN(n_0_0_402));
   AOI221_X1 i_0_0_409 (.A(n_0_0_404), .B1(B[17]), .B2(n_0_0_414), .C1(B[1]), 
      .C2(n_0_0_515), .ZN(n_0_0_403));
   INV_X1 i_0_0_410 (.A(n_0_0_405), .ZN(n_0_0_404));
   AOI22_X1 i_0_0_411 (.A1(n_0_0_594), .A2(n_0_0_556), .B1(B[9]), .B2(n_0_0_572), 
      .ZN(n_0_0_405));
   INV_X1 i_0_0_412 (.A(n_0_0_406), .ZN(n_27));
   AOI222_X1 i_0_0_413 (.A1(B[2]), .A2(n_48), .B1(n_0_0_600), .B2(n_0_0_411), 
      .C1(n_0_0_558), .C2(n_0_0_407), .ZN(n_0_0_406));
   AOI22_X1 i_0_0_414 (.A1(n_0_0_597), .A2(n_0_0_408), .B1(n_0_0_598), .B2(
      n_0_0_418), .ZN(n_0_0_407));
   AOI221_X1 i_0_0_415 (.A(n_0_0_409), .B1(B[10]), .B2(n_0_0_572), .C1(B[18]), 
      .C2(n_0_0_414), .ZN(n_0_0_408));
   OAI22_X1 i_0_0_416 (.A1(n_0_0_593), .A2(n_0_0_565), .B1(n_0_0_199), .B2(
      n_0_0_575), .ZN(n_0_0_409));
   OAI21_X1 i_0_0_417 (.A(n_0_0_410), .B1(n_0_0_202), .B2(n_0_0_617), .ZN(n_28));
   AOI22_X1 i_0_0_418 (.A1(n_0_0_600), .A2(n_0_0_417), .B1(n_0_0_558), .B2(
      n_0_0_411), .ZN(n_0_0_410));
   AOI22_X1 i_0_0_419 (.A1(n_0_0_597), .A2(n_0_0_412), .B1(n_0_0_598), .B2(
      n_0_0_555), .ZN(n_0_0_411));
   AOI221_X1 i_0_0_420 (.A(n_0_0_413), .B1(n_0_0_594), .B2(n_0_0_553), .C1(B[19]), 
      .C2(n_0_0_414), .ZN(n_0_0_412));
   OAI21_X1 i_0_0_421 (.A(n_0_0_415), .B1(n_0_0_202), .B2(n_0_0_575), .ZN(
      n_0_0_413));
   NOR3_X1 i_0_0_422 (.A1(n_0_0_592), .A2(n_0_0_590), .A3(n_0_0_594), .ZN(
      n_0_0_414));
   NAND2_X1 i_0_0_423 (.A1(B[11]), .A2(n_0_0_572), .ZN(n_0_0_415));
   INV_X1 i_0_0_424 (.A(n_0_0_416), .ZN(n_29));
   AOI222_X1 i_0_0_425 (.A1(n_0_0_558), .A2(n_0_0_417), .B1(B[4]), .B2(n_48), 
      .C1(n_0_0_600), .C2(n_0_0_551), .ZN(n_0_0_416));
   AOI22_X1 i_0_0_426 (.A1(n_0_0_597), .A2(n_0_0_418), .B1(n_0_0_598), .B2(
      n_0_0_561), .ZN(n_0_0_417));
   AOI222_X1 i_0_0_427 (.A1(B[16]), .A2(n_0_0_571), .B1(B[8]), .B2(n_0_0_576), 
      .C1(n_0_0_593), .C2(n_0_0_419), .ZN(n_0_0_418));
   OAI21_X1 i_0_0_428 (.A(n_0_0_420), .B1(n_0_0_201), .B2(n_0_0_577), .ZN(
      n_0_0_419));
   AOI22_X1 i_0_0_429 (.A1(B[12]), .A2(n_0_0_573), .B1(B[20]), .B2(n_0_0_566), 
      .ZN(n_0_0_420));
   INV_X1 i_0_0_430 (.A(n_0_0_426), .ZN(n_30));
   AOI222_X1 i_0_0_431 (.A1(n_0_0_600), .A2(n_0_0_432), .B1(B[6]), .B2(n_48), 
      .C1(n_0_0_558), .C2(n_0_0_560), .ZN(n_0_0_426));
   INV_X1 i_0_0_432 (.A(n_0_0_431), .ZN(n_31));
   AOI222_X1 i_0_0_433 (.A1(n_0_0_558), .A2(n_0_0_432), .B1(B[7]), .B2(n_48), 
      .C1(n_0_0_600), .C2(n_0_0_438), .ZN(n_0_0_431));
   AOI22_X1 i_0_0_434 (.A1(n_0_0_597), .A2(n_0_0_552), .B1(n_0_0_598), .B2(
      n_0_0_445), .ZN(n_0_0_432));
   INV_X1 i_0_0_435 (.A(n_0_0_437), .ZN(n_32));
   AOI222_X1 i_0_0_436 (.A1(n_0_0_558), .A2(n_0_0_438), .B1(B[8]), .B2(n_48), 
      .C1(n_0_0_600), .C2(n_0_0_444), .ZN(n_0_0_437));
   AOI22_X1 i_0_0_437 (.A1(n_0_0_597), .A2(n_0_0_568), .B1(n_0_0_598), .B2(
      n_0_0_448), .ZN(n_0_0_438));
   OAI21_X1 i_0_0_438 (.A(n_0_0_443), .B1(n_0_0_603), .B2(n_0_0_617), .ZN(n_33));
   AOI22_X1 i_0_0_439 (.A1(n_0_0_558), .A2(n_0_0_444), .B1(n_0_0_600), .B2(
      n_0_0_447), .ZN(n_0_0_443));
   AOI22_X1 i_0_0_440 (.A1(n_0_0_597), .A2(n_0_0_445), .B1(n_0_0_598), .B2(
      n_0_0_453), .ZN(n_0_0_444));
   AOI222_X1 i_0_0_441 (.A1(B[9]), .A2(n_0_0_515), .B1(n_0_0_479), .B2(n_0_0_573), 
      .C1(B[13]), .C2(n_0_0_576), .ZN(n_0_0_445));
   INV_X1 i_0_0_442 (.A(n_0_0_446), .ZN(n_34));
   AOI222_X1 i_0_0_443 (.A1(B[10]), .A2(n_48), .B1(n_0_0_600), .B2(n_0_0_452), 
      .C1(n_0_0_558), .C2(n_0_0_447), .ZN(n_0_0_446));
   AOI22_X1 i_0_0_444 (.A1(n_0_0_598), .A2(n_0_0_457), .B1(n_0_0_597), .B2(
      n_0_0_448), .ZN(n_0_0_447));
   INV_X1 i_0_0_445 (.A(n_0_0_449), .ZN(n_0_0_448));
   AOI22_X1 i_0_0_446 (.A1(n_0_0_594), .A2(n_0_0_466), .B1(n_0_0_593), .B2(
      n_0_0_567), .ZN(n_0_0_449));
   INV_X1 i_0_0_447 (.A(n_0_0_451), .ZN(n_35));
   AOI222_X1 i_0_0_448 (.A1(n_0_0_558), .A2(n_0_0_452), .B1(B[11]), .B2(n_48), 
      .C1(n_0_0_600), .C2(n_0_0_455), .ZN(n_0_0_451));
   AOI22_X1 i_0_0_449 (.A1(n_0_0_597), .A2(n_0_0_453), .B1(n_0_0_598), .B2(
      n_0_0_460), .ZN(n_0_0_452));
   AOI222_X1 i_0_0_450 (.A1(B[11]), .A2(n_0_0_515), .B1(n_0_0_491), .B2(
      n_0_0_573), .C1(B[15]), .C2(n_0_0_576), .ZN(n_0_0_453));
   OAI21_X1 i_0_0_451 (.A(n_0_0_454), .B1(n_0_0_606), .B2(n_0_0_617), .ZN(n_36));
   AOI22_X1 i_0_0_452 (.A1(n_0_0_600), .A2(n_0_0_459), .B1(n_0_0_558), .B2(
      n_0_0_455), .ZN(n_0_0_454));
   AOI22_X1 i_0_0_453 (.A1(n_0_0_597), .A2(n_0_0_457), .B1(n_0_0_465), .B2(
      n_0_0_456), .ZN(n_0_0_455));
   AOI21_X1 i_0_0_454 (.A(n_0_0_597), .B1(B[18]), .B2(n_0_0_576), .ZN(n_0_0_456));
   AOI222_X1 i_0_0_455 (.A1(B[16]), .A2(n_0_0_576), .B1(B[12]), .B2(n_0_0_515), 
      .C1(B[20]), .C2(n_0_0_572), .ZN(n_0_0_457));
   INV_X1 i_0_0_456 (.A(n_0_0_458), .ZN(n_37));
   AOI222_X1 i_0_0_457 (.A1(n_0_0_600), .A2(n_0_0_462), .B1(B[13]), .B2(n_48), 
      .C1(n_0_0_558), .C2(n_0_0_459), .ZN(n_0_0_458));
   AOI22_X1 i_0_0_458 (.A1(n_0_0_597), .A2(n_0_0_460), .B1(n_0_0_598), .B2(
      n_0_0_469), .ZN(n_0_0_459));
   AOI222_X1 i_0_0_459 (.A1(B[13]), .A2(n_0_0_515), .B1(B[21]), .B2(n_0_0_572), 
      .C1(B[17]), .C2(n_0_0_576), .ZN(n_0_0_460));
   INV_X1 i_0_0_460 (.A(n_0_0_461), .ZN(n_38));
   AOI222_X1 i_0_0_462 (.A1(B[14]), .A2(n_48), .B1(n_0_0_558), .B2(n_0_0_462), 
      .C1(n_0_0_600), .C2(n_0_0_468), .ZN(n_0_0_461));
   OAI21_X1 i_0_0_463 (.A(n_0_0_463), .B1(n_0_0_598), .B2(n_0_0_465), .ZN(
      n_0_0_462));
   AOI21_X1 i_0_0_464 (.A(n_0_0_464), .B1(n_0_0_486), .B2(n_0_0_576), .ZN(
      n_0_0_463));
   NOR3_X1 i_0_0_465 (.A1(n_0_0_608), .A2(n_0_0_597), .A3(n_0_0_575), .ZN(
      n_0_0_464));
   OR2_X1 i_0_0_466 (.A1(n_0_0_594), .A2(n_0_0_466), .ZN(n_0_0_465));
   AOI22_X1 i_0_0_467 (.A1(B[14]), .A2(n_0_0_589), .B1(B[22]), .B2(n_0_0_573), 
      .ZN(n_0_0_466));
   INV_X1 i_0_0_468 (.A(n_0_0_467), .ZN(n_39));
   AOI222_X1 i_0_0_469 (.A1(n_0_0_600), .A2(n_0_0_474), .B1(B[15]), .B2(n_48), 
      .C1(n_0_0_558), .C2(n_0_0_468), .ZN(n_0_0_467));
   OAI22_X1 i_0_0_470 (.A1(n_0_0_577), .A2(n_0_0_472), .B1(n_0_0_598), .B2(
      n_0_0_469), .ZN(n_0_0_468));
   AOI221_X1 i_0_0_471 (.A(n_0_0_572), .B1(B[19]), .B2(n_0_0_576), .C1(B[15]), 
      .C2(n_0_0_515), .ZN(n_0_0_469));
   NAND2_X1 i_0_0_472 (.A1(n_0_0_598), .A2(n_0_0_479), .ZN(n_0_0_472));
   INV_X1 i_0_0_473 (.A(n_0_0_473), .ZN(n_40));
   AOI222_X1 i_0_0_474 (.A1(n_0_0_558), .A2(n_0_0_474), .B1(B[16]), .B2(n_48), 
      .C1(n_0_0_600), .C2(n_0_0_478), .ZN(n_0_0_473));
   INV_X1 i_0_0_475 (.A(n_0_0_475), .ZN(n_0_0_474));
   AOI21_X1 i_0_0_476 (.A(n_0_0_476), .B1(n_0_0_498), .B2(n_0_0_576), .ZN(
      n_0_0_475));
   AOI221_X1 i_0_0_477 (.A(n_0_0_575), .B1(n_0_0_608), .B2(n_0_0_597), .C1(
      n_0_0_610), .C2(n_0_0_598), .ZN(n_0_0_476));
   INV_X1 i_0_0_478 (.A(n_0_0_477), .ZN(n_41));
   AOI222_X1 i_0_0_479 (.A1(n_0_0_558), .A2(n_0_0_478), .B1(B[17]), .B2(n_48), 
      .C1(n_0_0_600), .C2(n_0_0_482), .ZN(n_0_0_477));
   AOI221_X1 i_0_0_480 (.A(n_0_0_577), .B1(n_0_0_597), .B2(n_0_0_480), .C1(
      n_0_0_598), .C2(n_0_0_490), .ZN(n_0_0_478));
   INV_X1 i_0_0_481 (.A(n_0_0_480), .ZN(n_0_0_479));
   AOI22_X1 i_0_0_482 (.A1(B[17]), .A2(n_0_0_593), .B1(B[21]), .B2(n_0_0_594), 
      .ZN(n_0_0_480));
   INV_X1 i_0_0_483 (.A(n_0_0_481), .ZN(n_42));
   AOI222_X1 i_0_0_484 (.A1(n_0_0_558), .A2(n_0_0_482), .B1(B[18]), .B2(n_48), 
      .C1(n_0_0_600), .C2(n_0_0_488), .ZN(n_0_0_481));
   OAI21_X1 i_0_0_485 (.A(n_0_0_485), .B1(n_0_0_613), .B2(n_0_0_483), .ZN(
      n_0_0_482));
   NAND2_X1 i_0_0_486 (.A1(n_0_0_597), .A2(n_0_0_576), .ZN(n_0_0_483));
   NAND2_X1 i_0_0_487 (.A1(n_0_0_515), .A2(n_0_0_486), .ZN(n_0_0_485));
   OAI22_X1 i_0_0_488 (.A1(n_0_0_610), .A2(n_0_0_598), .B1(n_0_0_612), .B2(
      n_0_0_597), .ZN(n_0_0_486));
   INV_X1 i_0_0_489 (.A(n_0_0_487), .ZN(n_43));
   AOI221_X1 i_0_0_490 (.A(n_0_0_494), .B1(n_0_0_558), .B2(n_0_0_488), .C1(B[19]), 
      .C2(n_48), .ZN(n_0_0_487));
   AOI211_X1 i_0_0_491 (.A(n_0_0_489), .B(n_0_0_577), .C1(n_0_0_597), .C2(
      n_0_0_490), .ZN(n_0_0_488));
   AOI21_X1 i_0_0_492 (.A(n_0_0_597), .B1(B[21]), .B2(n_0_0_593), .ZN(n_0_0_489));
   INV_X1 i_0_0_493 (.A(n_0_0_491), .ZN(n_0_0_490));
   NAND2_X1 i_0_0_494 (.A1(n_0_0_611), .A2(n_0_0_593), .ZN(n_0_0_491));
   AND3_X1 i_0_0_495 (.A1(n_0_0_515), .A2(n_0_0_498), .A3(n_0_0_600), .ZN(
      n_0_0_494));
   INV_X1 i_0_0_496 (.A(n_0_0_496), .ZN(n_44));
   AOI22_X1 i_0_0_497 (.A1(B[20]), .A2(n_48), .B1(n_0_0_601), .B2(n_0_0_497), 
      .ZN(n_0_0_496));
   AOI211_X1 i_0_0_498 (.A(n_0_0_500), .B(n_0_0_575), .C1(n_0_0_540), .C2(
      n_0_0_499), .ZN(n_0_0_497));
   INV_X1 i_0_0_499 (.A(n_0_0_499), .ZN(n_0_0_498));
   AOI22_X1 i_0_0_500 (.A1(B[22]), .A2(n_0_0_598), .B1(B[20]), .B2(n_0_0_597), 
      .ZN(n_0_0_499));
   NOR3_X1 i_0_0_603 (.A1(B[21]), .A2(n_0_0_598), .A3(n_0_0_540), .ZN(n_0_0_500));
   INV_X1 i_0_0_501 (.A(n_0_0_501), .ZN(n_45));
   AOI22_X1 i_0_0_502 (.A1(B[21]), .A2(n_48), .B1(n_0_0_601), .B2(n_0_0_502), 
      .ZN(n_0_0_501));
   AOI211_X1 i_0_0_503 (.A(n_0_0_470), .B(n_0_0_575), .C1(n_0_0_613), .C2(
      n_0_0_539), .ZN(n_0_0_502));
   AOI21_X1 i_0_0_504 (.A(n_0_0_532), .B1(n_0_0_617), .B2(n_0_0_504), .ZN(n_46));
   NAND3_X1 i_0_0_505 (.A1(n_0_0_602), .A2(n_0_0_597), .A3(n_0_0_515), .ZN(
      n_0_0_504));
   INV_X1 i_0_0_506 (.A(n_0_0_575), .ZN(n_0_0_515));
   AOI22_X1 i_0_0_507 (.A1(B[24]), .A2(n_0_0_96), .B1(B[23]), .B2(n_0_0_547), 
      .ZN(n_0_0_95));
   AOI21_X1 i_0_0_508 (.A(B[22]), .B1(n_0_0_617), .B2(n_0_0_539), .ZN(n_0_0_532));
   INV_X1 i_0_0_509 (.A(n_0_0_538), .ZN(exp_Sum[7]));
   INV_X1 i_0_0_510 (.A(n_0_0_6), .ZN(n_0_0_563));
   INV_X1 i_0_0_511 (.A(n_0_28), .ZN(n_0_0_564));
   INV_X1 i_0_0_685 (.A(A[12]), .ZN(n_0_0_578));
   INV_X1 i_0_0_512 (.A(A[13]), .ZN(n_0_0_579));
   INV_X1 i_0_0_687 (.A(A[14]), .ZN(n_0_0_580));
   INV_X1 i_0_0_688 (.A(A[15]), .ZN(n_0_0_581));
   INV_X1 i_0_0_689 (.A(A[16]), .ZN(n_0_0_582));
   INV_X1 i_0_0_690 (.A(A[17]), .ZN(n_0_0_583));
   INV_X1 i_0_0_691 (.A(A[18]), .ZN(n_0_0_584));
   INV_X1 i_0_0_692 (.A(A[19]), .ZN(n_0_0_585));
   INV_X1 i_0_0_513 (.A(A[20]), .ZN(n_0_0_586));
   INV_X1 i_0_0_514 (.A(A[21]), .ZN(n_0_0_587));
   INV_X1 i_0_0_515 (.A(A[22]), .ZN(n_0_0_588));
   INV_X1 i_0_0_516 (.A(A[24]), .ZN(n_0_0_96));
   INV_X1 i_0_0_517 (.A(B[9]), .ZN(n_0_0_603));
   INV_X1 i_0_0_711 (.A(B[10]), .ZN(n_0_0_604));
   INV_X1 i_0_0_712 (.A(B[11]), .ZN(n_0_0_605));
   INV_X1 i_0_0_518 (.A(B[12]), .ZN(n_0_0_606));
   INV_X1 i_0_0_714 (.A(B[13]), .ZN(n_0_0_607));
   INV_X1 i_0_0_519 (.A(B[16]), .ZN(n_0_0_608));
   INV_X1 i_0_0_716 (.A(B[17]), .ZN(n_0_0_609));
   INV_X1 i_0_0_520 (.A(B[18]), .ZN(n_0_0_610));
   INV_X1 i_0_0_521 (.A(B[19]), .ZN(n_0_0_611));
   INV_X1 i_0_0_522 (.A(B[20]), .ZN(n_0_0_612));
   INV_X1 i_0_0_523 (.A(B[22]), .ZN(n_0_0_613));
   INV_X1 i_0_0_524 (.A(B[25]), .ZN(n_0_0_99));
   INV_X1 i_0_0_525 (.A(B[31]), .ZN(n_0_0_94));
   OAI22_X1 i_0_0_526 (.A1(n_0_1), .A2(n_0_0_110), .B1(n_0_0_125), .B2(n_0_0_101), 
      .ZN(n_0_0_100));
   AOI22_X1 i_0_0_527 (.A1(n_0_0_126), .A2(n_0_0_102), .B1(n_0_2), .B2(n_0_0_109), 
      .ZN(n_0_0_101));
   AOI222_X1 i_0_0_528 (.A1(n_9), .A2(n_0_0_120), .B1(n_1), .B2(n_0_0_122), 
      .C1(n_17), .C2(n_0_0_114), .ZN(n_0_0_102));
   AOI22_X1 i_0_0_529 (.A1(n_13), .A2(n_0_0_114), .B1(n_5), .B2(n_0_0_120), 
      .ZN(n_0_0_109));
   OAI21_X1 i_0_0_530 (.A(n_0_0_111), .B1(n_0_0_126), .B2(n_0_0_112), .ZN(
      n_0_0_110));
   AOI222_X1 i_0_0_531 (.A1(n_19), .A2(n_0_0_113), .B1(n_11), .B2(n_0_0_119), 
      .C1(n_3), .C2(n_0_0_121), .ZN(n_0_0_111));
   AOI22_X1 i_0_0_532 (.A1(n_15), .A2(n_0_0_114), .B1(n_7), .B2(n_0_0_120), 
      .ZN(n_0_0_112));
   NOR3_X1 i_0_0_533 (.A1(n_0_4), .A2(n_0_3), .A3(n_0_2), .ZN(n_0_0_113));
   NOR2_X1 i_0_0_534 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_0_114));
   NOR3_X1 i_0_0_535 (.A1(n_0_4), .A2(n_0_0_128), .A3(n_0_2), .ZN(n_0_0_119));
   NOR2_X1 i_0_0_536 (.A1(n_0_4), .A2(n_0_0_128), .ZN(n_0_0_120));
   NOR3_X1 i_0_0_537 (.A1(n_0_0_129), .A2(n_0_3), .A3(n_0_2), .ZN(n_0_0_121));
   NOR2_X1 i_0_0_538 (.A1(n_0_0_129), .A2(n_0_3), .ZN(n_0_0_122));
   INV_X1 i_0_0_539 (.A(n_0_1), .ZN(n_0_0_125));
   INV_X1 i_0_0_540 (.A(n_0_2), .ZN(n_0_0_126));
   INV_X1 i_0_0_541 (.A(n_0_3), .ZN(n_0_0_128));
   INV_X1 i_0_0_542 (.A(n_0_4), .ZN(n_0_0_129));
   OAI21_X1 i_0_0_543 (.A(n_0_0_131), .B1(n_0_1), .B2(n_0_0_132), .ZN(n_0_0_130));
   NAND2_X1 i_0_0_544 (.A1(n_0_1), .A2(n_0_0_195), .ZN(n_0_0_131));
   INV_X1 i_0_0_545 (.A(n_0_0_192), .ZN(n_0_0_132));
   OAI21_X1 i_0_0_546 (.A(n_0_0_193), .B1(n_0_0_126), .B2(n_0_0_194), .ZN(
      n_0_0_192));
   AOI222_X1 i_0_0_547 (.A1(n_20), .A2(n_0_0_113), .B1(n_12), .B2(n_0_0_119), 
      .C1(n_4), .C2(n_0_0_121), .ZN(n_0_0_193));
   AOI222_X1 i_0_0_548 (.A1(n_16), .A2(n_0_0_114), .B1(n_0), .B2(n_0_0_122), 
      .C1(n_8), .C2(n_0_0_120), .ZN(n_0_0_194));
   OAI22_X1 i_0_0_549 (.A1(n_0_2), .A2(n_0_0_197), .B1(n_0_0_126), .B2(n_0_0_196), 
      .ZN(n_0_0_195));
   AOI22_X1 i_0_0_550 (.A1(n_14), .A2(n_0_0_114), .B1(n_6), .B2(n_0_0_120), 
      .ZN(n_0_0_196));
   AOI222_X1 i_0_0_551 (.A1(n_18), .A2(n_0_0_114), .B1(n_2), .B2(n_0_0_122), 
      .C1(n_10), .C2(n_0_0_120), .ZN(n_0_0_197));
   INV_X1 i_0_0_552 (.A(A[1]), .ZN(n_0_0_198));
   INV_X1 i_0_0_553 (.A(B[2]), .ZN(n_0_0_199));
   INV_X1 i_0_0_554 (.A(B[1]), .ZN(n_0_0_200));
   INV_X1 i_0_0_555 (.A(B[4]), .ZN(n_0_0_201));
   INV_X1 i_0_0_556 (.A(B[3]), .ZN(n_0_0_202));
   INV_X1 i_0_0_557 (.A(A[4]), .ZN(n_0_0_306));
   INV_X1 i_0_0_558 (.A(A[5]), .ZN(n_0_0_307));
   INV_X1 i_0_0_559 (.A(B[5]), .ZN(n_0_0_308));
   INV_X1 i_0_0_560 (.A(A[6]), .ZN(n_0_0_309));
   INV_X1 i_0_0_561 (.A(A[7]), .ZN(n_0_0_310));
   INV_X1 i_0_0_562 (.A(B[7]), .ZN(n_0_0_312));
   INV_X1 i_0_0_563 (.A(A[8]), .ZN(n_0_0_313));
   INV_X1 i_0_0_564 (.A(B[8]), .ZN(n_0_0_314));
   INV_X1 i_0_0_565 (.A(A[0]), .ZN(n_0_0_315));
   OAI22_X1 i_0_0_566 (.A1(n_0_0_315), .A2(B[0]), .B1(n_0_0_198), .B2(B[1]), 
      .ZN(n_0_0_316));
   OAI221_X1 i_0_0_567 (.A(n_0_0_316), .B1(n_0_0_199), .B2(A[2]), .C1(n_0_0_200), 
      .C2(A[1]), .ZN(n_0_0_319));
   INV_X1 i_0_0_568 (.A(A[3]), .ZN(n_0_0_323));
   INV_X1 i_0_0_569 (.A(A[2]), .ZN(n_0_0_324));
   OAI221_X1 i_0_0_570 (.A(n_0_0_319), .B1(B[3]), .B2(n_0_0_323), .C1(n_0_0_324), 
      .C2(B[2]), .ZN(n_0_0_325));
   OAI221_X1 i_0_0_571 (.A(n_0_0_325), .B1(A[4]), .B2(n_0_0_201), .C1(n_0_0_202), 
      .C2(A[3]), .ZN(n_0_0_326));
   OAI221_X1 i_0_0_572 (.A(n_0_0_326), .B1(n_0_0_306), .B2(B[4]), .C1(B[5]), 
      .C2(n_0_0_307), .ZN(n_0_0_327));
   INV_X1 i_0_0_573 (.A(B[6]), .ZN(n_0_0_333));
   OAI221_X1 i_0_0_574 (.A(n_0_0_327), .B1(A[6]), .B2(n_0_0_333), .C1(n_0_0_308), 
      .C2(A[5]), .ZN(n_0_0_345));
   OAI221_X1 i_0_0_575 (.A(n_0_0_345), .B1(n_0_0_309), .B2(B[6]), .C1(B[7]), 
      .C2(n_0_0_310), .ZN(n_0_0_352));
   NAND2_X1 i_0_0_576 (.A1(n_0_0_310), .A2(B[7]), .ZN(n_0_0_353));
   AOI22_X1 i_0_0_577 (.A1(n_0_0_352), .A2(n_0_0_353), .B1(n_0_0_314), .B2(A[8]), 
      .ZN(n_0_0_354));
   INV_X1 i_0_0_578 (.A(A[9]), .ZN(n_0_0_361));
   AOI221_X1 i_0_0_579 (.A(n_0_0_354), .B1(B[8]), .B2(n_0_0_313), .C1(B[9]), 
      .C2(n_0_0_361), .ZN(n_0_0_362));
   INV_X1 i_0_0_580 (.A(n_0_0_366), .ZN(n_0_36));
   AOI222_X1 i_0_0_581 (.A1(n_0_0_484), .A2(n_0_0_391), .B1(A[7]), .B2(n_0_52), 
      .C1(n_0_0_390), .C2(n_0_0_369), .ZN(n_0_0_366));
   AOI22_X1 i_0_0_582 (.A1(n_0_0_470), .A2(n_0_0_374), .B1(n_0_0_450), .B2(
      n_0_0_385), .ZN(n_0_0_369));
   AOI221_X1 i_0_0_583 (.A(n_0_0_375), .B1(A[16]), .B2(n_0_0_388), .C1(A[20]), 
      .C2(n_0_0_389), .ZN(n_0_0_374));
   OAI21_X1 i_0_0_584 (.A(n_0_0_383), .B1(n_0_0_313), .B2(n_0_0_421), .ZN(
      n_0_0_375));
   NAND2_X1 i_0_0_585 (.A1(A[12]), .A2(n_0_0_394), .ZN(n_0_0_383));
   INV_X1 i_0_0_586 (.A(n_0_0_385), .ZN(n_0_0_384));
   AOI221_X1 i_0_0_587 (.A(n_0_0_386), .B1(A[22]), .B2(n_0_0_389), .C1(A[10]), 
      .C2(n_0_0_422), .ZN(n_0_0_385));
   INV_X1 i_0_0_588 (.A(n_0_0_387), .ZN(n_0_0_386));
   AOI22_X1 i_0_0_589 (.A1(A[18]), .A2(n_0_0_388), .B1(A[14]), .B2(n_0_0_394), 
      .ZN(n_0_0_387));
   NOR2_X1 i_0_0_590 (.A1(n_0_0_441), .A2(n_0_0_434), .ZN(n_0_0_388));
   NOR2_X1 i_0_0_591 (.A1(n_0_0_442), .A2(n_0_0_434), .ZN(n_0_0_389));
   NOR2_X1 i_0_0_592 (.A1(n_0_0_540), .A2(n_0_0_493), .ZN(n_0_0_390));
   OAI22_X1 i_0_0_593 (.A1(n_0_0_470), .A2(n_0_0_392), .B1(n_0_0_450), .B2(
      n_0_0_423), .ZN(n_0_0_391));
   AOI221_X1 i_0_0_594 (.A(n_0_0_393), .B1(A[9]), .B2(n_0_0_422), .C1(A[13]), 
      .C2(n_0_0_394), .ZN(n_0_0_392));
   NOR2_X1 i_0_0_595 (.A1(n_0_0_434), .A2(n_0_0_395), .ZN(n_0_0_393));
   NOR2_X1 i_0_0_596 (.A1(n_0_0_442), .A2(n_0_0_430), .ZN(n_0_0_394));
   OAI22_X1 i_0_0_597 (.A1(A[21]), .A2(n_0_0_442), .B1(A[17]), .B2(n_0_0_441), 
      .ZN(n_0_0_395));
   INV_X1 i_0_0_598 (.A(n_0_0_422), .ZN(n_0_0_421));
   NOR2_X1 i_0_0_599 (.A1(n_0_0_441), .A2(n_0_0_430), .ZN(n_0_0_422));
   OAI22_X1 i_0_0_600 (.A1(n_0_0_441), .A2(n_0_0_424), .B1(n_0_0_442), .B2(
      n_0_0_427), .ZN(n_0_0_423));
   AOI22_X1 i_0_0_601 (.A1(n_0_0_439), .A2(n_0_0_425), .B1(n_0_0_310), .B2(
      n_0_0_429), .ZN(n_0_0_424));
   NAND2_X1 i_0_0_602 (.A1(A[15]), .A2(n_0_0_435), .ZN(n_0_0_425));
   INV_X1 i_0_0_604 (.A(n_0_0_428), .ZN(n_0_0_427));
   AOI22_X1 i_0_0_605 (.A1(A[11]), .A2(n_0_0_429), .B1(A[19]), .B2(n_0_0_433), 
      .ZN(n_0_0_428));
   INV_X1 i_0_0_606 (.A(n_0_0_430), .ZN(n_0_0_429));
   NAND2_X1 i_0_0_607 (.A1(n_0_0_440), .A2(n_0_0_435), .ZN(n_0_0_430));
   INV_X1 i_0_0_608 (.A(n_0_0_434), .ZN(n_0_0_433));
   NAND2_X1 i_0_0_609 (.A1(n_0_0_439), .A2(n_0_0_435), .ZN(n_0_0_434));
   XOR2_X1 i_0_0_610 (.A(n_0_0_507), .B(n_0_0_436), .Z(n_0_0_435));
   OAI21_X1 i_0_0_611 (.A(n_0_0_522), .B1(A[27]), .B2(n_0_0_543), .ZN(n_0_0_436));
   INV_X1 i_0_0_612 (.A(n_0_0_440), .ZN(n_0_0_439));
   XOR2_X1 i_0_0_613 (.A(n_0_0_526), .B(n_0_0_508), .Z(n_0_0_440));
   INV_X1 i_0_0_614 (.A(n_0_0_442), .ZN(n_0_0_441));
   XOR2_X1 i_0_0_615 (.A(n_0_0_512), .B(n_0_0_509), .Z(n_0_0_442));
   INV_X1 i_0_0_616 (.A(n_0_0_470), .ZN(n_0_0_450));
   XOR2_X1 i_0_0_617 (.A(n_0_0_541), .B(n_0_0_511), .Z(n_0_0_470));
   INV_X1 i_0_0_618 (.A(n_0_0_484), .ZN(n_0_0_471));
   NOR2_X1 i_0_0_619 (.A1(n_0_0_539), .A2(n_0_0_493), .ZN(n_0_0_484));
   INV_X1 i_0_0_620 (.A(n_0_0_493), .ZN(n_0_0_492));
   OAI221_X1 i_0_0_621 (.A(n_0_0_516), .B1(n_0_0_519), .B2(n_0_0_506), .C1(
      n_0_0_505), .C2(n_0_0_495), .ZN(n_0_0_493));
   OAI33_X1 i_0_0_622 (.A1(n_0_0_549), .A2(B[28]), .A3(n_0_0_503), .B1(A[28]), 
      .B2(n_0_0_544), .B3(n_0_0_531), .ZN(n_0_0_495));
   AOI22_X1 i_0_0_623 (.A1(A[29]), .A2(n_0_0_545), .B1(n_0_0_536), .B2(n_0_0_534), 
      .ZN(n_0_0_503));
   INV_X1 i_0_0_624 (.A(n_0_0_506), .ZN(n_0_0_505));
   AOI21_X1 i_0_0_625 (.A(n_0_0_521), .B1(n_0_0_522), .B2(n_0_0_507), .ZN(
      n_0_0_506));
   AOI22_X1 i_0_0_626 (.A1(A[26]), .A2(n_0_0_542), .B1(n_0_0_526), .B2(n_0_0_508), 
      .ZN(n_0_0_507));
   OAI22_X1 i_0_0_627 (.A1(n_0_0_548), .A2(B[25]), .B1(n_0_0_512), .B2(n_0_0_509), 
      .ZN(n_0_0_508));
   AOI21_X1 i_0_0_628 (.A(n_0_0_514), .B1(n_0_0_541), .B2(n_0_0_511), .ZN(
      n_0_0_509));
   INV_X1 i_0_0_629 (.A(n_0_0_511), .ZN(n_0_0_510));
   AOI21_X1 i_0_0_630 (.A(n_0_0_514), .B1(B[24]), .B2(n_0_0_96), .ZN(n_0_0_511));
   INV_X1 i_0_0_631 (.A(n_0_0_513), .ZN(n_0_0_512));
   OAI22_X1 i_0_0_632 (.A1(A[25]), .A2(B[25]), .B1(n_0_0_548), .B2(n_0_0_99), 
      .ZN(n_0_0_513));
   NOR2_X1 i_0_0_633 (.A1(B[24]), .A2(n_0_0_96), .ZN(n_0_0_514));
   INV_X1 i_0_0_634 (.A(n_0_52), .ZN(n_0_0_516));
   NAND2_X1 i_0_0_635 (.A1(n_0_0_527), .A2(n_0_0_517), .ZN(n_0_52));
   NAND3_X1 i_0_0_636 (.A1(n_0_0_527), .A2(n_0_0_520), .A3(n_0_0_519), .ZN(
      n_0_0_517));
   INV_X1 i_0_0_637 (.A(n_0_0_519), .ZN(n_0_0_518));
   AOI211_X1 i_0_0_638 (.A(n_0_0_529), .B(n_0_0_534), .C1(n_0_0_549), .C2(B[28]), 
      .ZN(n_0_0_519));
   OAI21_X1 i_0_0_639 (.A(n_0_0_522), .B1(n_0_0_523), .B2(n_0_0_521), .ZN(
      n_0_0_520));
   NOR2_X1 i_0_0_640 (.A1(A[27]), .A2(n_0_0_543), .ZN(n_0_0_521));
   NAND2_X1 i_0_0_641 (.A1(A[27]), .A2(n_0_0_543), .ZN(n_0_0_522));
   OAI21_X1 i_0_0_642 (.A(n_0_0_524), .B1(A[26]), .B2(n_0_0_542), .ZN(n_0_0_523));
   NAND2_X1 i_0_0_643 (.A1(n_0_0_526), .A2(n_0_0_525), .ZN(n_0_0_524));
   OAI21_X1 i_0_0_644 (.A(n_0_0_595), .B1(A[25]), .B2(n_0_0_99), .ZN(n_0_0_525));
   XOR2_X1 i_0_0_645 (.A(A[26]), .B(n_0_0_542), .Z(n_0_0_526));
   NOR2_X1 i_0_0_646 (.A1(n_0_0_530), .A2(n_0_0_528), .ZN(n_0_0_527));
   NOR2_X1 i_0_0_647 (.A1(n_0_0_535), .A2(n_0_0_529), .ZN(n_0_0_528));
   NOR2_X1 i_0_0_648 (.A1(A[30]), .A2(n_0_0_546), .ZN(n_0_0_529));
   NOR3_X1 i_0_0_649 (.A1(n_0_0_549), .A2(B[28]), .A3(n_0_0_531), .ZN(n_0_0_530));
   NAND2_X1 i_0_0_650 (.A1(n_0_0_535), .A2(n_0_0_533), .ZN(n_0_0_531));
   INV_X1 i_0_0_651 (.A(n_0_0_534), .ZN(n_0_0_533));
   NOR2_X1 i_0_0_652 (.A1(A[29]), .A2(n_0_0_545), .ZN(n_0_0_534));
   AOI21_X1 i_0_0_653 (.A(n_0_0_537), .B1(A[29]), .B2(n_0_0_545), .ZN(n_0_0_535));
   INV_X1 i_0_0_654 (.A(n_0_0_537), .ZN(n_0_0_536));
   AOI21_X1 i_0_0_655 (.A(n_0_0_538), .B1(A[30]), .B2(B[30]), .ZN(n_0_0_537));
   NOR2_X1 i_0_0_656 (.A1(A[30]), .A2(B[30]), .ZN(n_0_0_538));
   INV_X1 i_0_0_657 (.A(n_0_0_540), .ZN(n_0_0_539));
   AOI21_X1 i_0_0_658 (.A(n_0_0_541), .B1(n_0_0_547), .B2(B[23]), .ZN(n_0_0_540));
   NOR2_X1 i_0_0_659 (.A1(n_0_0_547), .A2(B[23]), .ZN(n_0_0_541));
   INV_X1 i_0_0_660 (.A(B[26]), .ZN(n_0_0_542));
   INV_X1 i_0_0_661 (.A(B[27]), .ZN(n_0_0_543));
   INV_X1 i_0_0_662 (.A(B[28]), .ZN(n_0_0_544));
   INV_X1 i_0_0_663 (.A(B[29]), .ZN(n_0_0_545));
   INV_X1 i_0_0_664 (.A(B[30]), .ZN(n_0_0_546));
   INV_X1 i_0_0_665 (.A(A[23]), .ZN(n_0_0_547));
   INV_X1 i_0_0_666 (.A(A[25]), .ZN(n_0_0_548));
   INV_X1 i_0_0_667 (.A(A[28]), .ZN(n_0_0_549));
   INV_X1 i_0_0_668 (.A(n_0_0_550), .ZN(n_47));
   AOI222_X1 i_0_0_669 (.A1(n_0_0_600), .A2(n_0_0_560), .B1(B[5]), .B2(n_48), 
      .C1(n_0_0_558), .C2(n_0_0_551), .ZN(n_0_0_550));
   OAI22_X1 i_0_0_670 (.A1(n_0_0_597), .A2(n_0_0_552), .B1(n_0_0_598), .B2(
      n_0_0_555), .ZN(n_0_0_551));
   AOI222_X1 i_0_0_671 (.A1(n_0_0_593), .A2(n_0_0_553), .B1(B[11]), .B2(
      n_0_0_576), .C1(B[19]), .C2(n_0_0_571), .ZN(n_0_0_552));
   AOI22_X1 i_0_0_672 (.A1(n_0_0_592), .A2(n_0_0_554), .B1(n_0_0_312), .B2(
      n_0_0_589), .ZN(n_0_0_553));
   NAND2_X1 i_0_0_673 (.A1(B[15]), .A2(n_0_0_590), .ZN(n_0_0_554));
   AOI222_X1 i_0_0_674 (.A1(B[9]), .A2(n_0_0_576), .B1(B[17]), .B2(n_0_0_571), 
      .C1(n_0_0_593), .C2(n_0_0_556), .ZN(n_0_0_555));
   OAI21_X1 i_0_0_675 (.A(n_0_0_557), .B1(n_0_0_308), .B2(n_0_0_577), .ZN(
      n_0_0_556));
   AOI22_X1 i_0_0_676 (.A1(B[21]), .A2(n_0_0_566), .B1(B[13]), .B2(n_0_0_573), 
      .ZN(n_0_0_557));
   INV_X1 i_0_0_677 (.A(n_0_0_559), .ZN(n_0_0_558));
   NAND2_X1 i_0_0_678 (.A1(n_0_0_540), .A2(n_0_0_601), .ZN(n_0_0_559));
   OAI22_X1 i_0_0_679 (.A1(n_0_0_598), .A2(n_0_0_561), .B1(n_0_0_597), .B2(
      n_0_0_568), .ZN(n_0_0_560));
   INV_X1 i_0_0_680 (.A(n_0_0_562), .ZN(n_0_0_561));
   OAI22_X1 i_0_0_681 (.A1(n_0_0_594), .A2(n_0_0_565), .B1(n_0_0_593), .B2(
      n_0_0_567), .ZN(n_0_0_562));
   AOI222_X1 i_0_0_682 (.A1(B[22]), .A2(n_0_0_566), .B1(B[6]), .B2(n_0_0_589), 
      .C1(B[14]), .C2(n_0_0_573), .ZN(n_0_0_565));
   NOR2_X1 i_0_0_683 (.A1(n_0_0_592), .A2(n_0_0_590), .ZN(n_0_0_566));
   AOI22_X1 i_0_0_684 (.A1(B[10]), .A2(n_0_0_589), .B1(B[18]), .B2(n_0_0_573), 
      .ZN(n_0_0_567));
   AOI221_X1 i_0_0_686 (.A(n_0_0_569), .B1(B[16]), .B2(n_0_0_572), .C1(B[20]), 
      .C2(n_0_0_571), .ZN(n_0_0_568));
   OAI21_X1 i_0_0_693 (.A(n_0_0_570), .B1(n_0_0_314), .B2(n_0_0_575), .ZN(
      n_0_0_569));
   NAND2_X1 i_0_0_694 (.A1(B[12]), .A2(n_0_0_576), .ZN(n_0_0_570));
   NOR2_X1 i_0_0_695 (.A1(n_0_0_593), .A2(n_0_0_574), .ZN(n_0_0_571));
   NOR2_X1 i_0_0_696 (.A1(n_0_0_594), .A2(n_0_0_574), .ZN(n_0_0_572));
   INV_X1 i_0_0_697 (.A(n_0_0_574), .ZN(n_0_0_573));
   NAND2_X1 i_0_0_698 (.A1(n_0_0_592), .A2(n_0_0_590), .ZN(n_0_0_574));
   NAND2_X1 i_0_0_699 (.A1(n_0_0_593), .A2(n_0_0_589), .ZN(n_0_0_575));
   NOR2_X1 i_0_0_700 (.A1(n_0_0_593), .A2(n_0_0_577), .ZN(n_0_0_576));
   INV_X1 i_0_0_701 (.A(n_0_0_589), .ZN(n_0_0_577));
   NOR2_X1 i_0_0_702 (.A1(n_0_0_592), .A2(n_0_0_591), .ZN(n_0_0_589));
   INV_X1 i_0_0_703 (.A(n_0_0_591), .ZN(n_0_0_590));
   XOR2_X1 i_0_0_704 (.A(n_0_0_523), .B(n_0_0_436), .Z(n_0_0_591));
   OAI21_X1 i_0_0_705 (.A(n_0_0_524), .B1(n_0_0_526), .B2(n_0_0_525), .ZN(
      n_0_0_592));
   INV_X1 i_0_0_706 (.A(n_0_0_594), .ZN(n_0_0_593));
   OAI21_X1 i_0_0_707 (.A(n_0_0_595), .B1(n_0_0_513), .B2(n_0_0_596), .ZN(
      n_0_0_594));
   NAND2_X1 i_0_0_708 (.A1(n_0_0_513), .A2(n_0_0_596), .ZN(n_0_0_595));
   NOR2_X1 i_0_0_709 (.A1(n_0_0_514), .A2(n_0_0_95), .ZN(n_0_0_596));
   INV_X1 i_0_0_710 (.A(n_0_0_598), .ZN(n_0_0_597));
   OAI21_X1 i_0_0_713 (.A(n_0_0_599), .B1(n_0_0_540), .B2(n_0_0_450), .ZN(
      n_0_0_598));
   NAND2_X1 i_0_0_715 (.A1(n_0_0_510), .A2(n_0_0_540), .ZN(n_0_0_599));
   AND2_X1 i_0_0_717 (.A1(n_0_0_539), .A2(n_0_0_601), .ZN(n_0_0_600));
   AND2_X1 i_0_0_718 (.A1(n_0_0_617), .A2(n_0_0_602), .ZN(n_0_0_601));
   OAI21_X1 i_0_0_719 (.A(n_0_0_517), .B1(n_0_0_520), .B2(n_0_0_614), .ZN(
      n_0_0_602));
   AOI21_X1 i_0_0_720 (.A(n_0_0_530), .B1(n_0_0_616), .B2(n_0_0_615), .ZN(
      n_0_0_614));
   NOR3_X1 i_0_0_721 (.A1(n_0_0_535), .A2(A[28]), .A3(n_0_0_544), .ZN(n_0_0_615));
   NAND2_X1 i_0_0_722 (.A1(n_0_0_537), .A2(n_0_0_533), .ZN(n_0_0_616));
   INV_X1 i_0_0_723 (.A(n_0_0_617), .ZN(n_48));
   OAI21_X1 i_0_0_724 (.A(n_0_0_527), .B1(n_0_0_518), .B2(n_0_0_505), .ZN(
      n_0_0_617));
endmodule
